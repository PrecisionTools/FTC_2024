.subckt AD3552R_INL code INL
E1 INL 0 code 0 table = (0,0.000000), (1,-0.026886), (2,0.234685), (3,0.117687), (4,0.037389), (5,-0.148356), (6,0.223295), (7,0.079823), (8,0.101246), (9,-0.050122), (10,0.386562), (11,0.218006), (12,0.181834), (13,-0.019703), (14,0.256263), (15,0.131376), (16,0.022738), (17,-0.130020), (18,0.205864), (19,0.054032), (20,-0.017443), (21,-0.192969), (22,0.173579), (23,0.004559), (24,0.062675), (25,-0.088229), (26,0.316865), (27,0.166430), (28,0.123752), (29,-0.046664), (30,0.184249), (31,0.038918), (32,-0.024662), (33,-0.190425), (34,0.352157), (35,0.209618), (36,0.131173), (37,0.007212), (38,0.392332), (39,0.224245), (40,0.069158), (41,-0.047840), (42,0.361437), (43,0.153401), (44,0.126515), (45,-0.029963), (46,0.237644), (47,0.084886), (48,0.029666), (49,-0.113806), (50,0.400912), (51,0.281127), (52,0.205006), (53,0.055961), (54,0.406247), (55,0.239550), (56,0.055202), (57,-0.130073), (58,0.301965), (59,0.148274), (60,0.084232), (61,-0.061564), (62,0.197214), (63,0.059315), (64,-0.023306), (65,-0.188613), (66,0.370700), (67,0.219332), (68,0.175258), (69,0.029926), (70,0.404833), (71,0.224668), (72,0.016162), (73,-0.160284), (74,0.271748), (75,0.105984), (76,0.057734), (77,-0.115469), (78,0.156321), (79,0.020745), (80,-0.036335), (81,-0.203495), (82,0.329337), (83,0.214199), (84,0.126932), (85,-0.024436), (86,0.336996), (87,0.198170), (88,0.002676), (89,-0.125931), (90,0.261512), (91,0.134758), (92,0.027053), (93,-0.105267), (94,0.152121), (95,-0.027118), (96,-0.063760), (97,-0.199799), (98,0.324674), (99,0.176092), (100,0.116226), (101,-0.058366), (102,0.330009), (103,0.144734), (104,-0.077704), (105,0.208945), (106,0.232691), (107,0.053922), (108,0.006134), (109,-0.184250), (110,0.073601), (111,-0.031788), (112,-0.107440), (113,0.134150), (114,0.293993), (115,0.153777), (116,0.090198), (117,0.039624), (118,0.326736), (119,0.130315), (120,0.024000), (121,-0.100894), (122,0.289342), (123,0.133327), (124,0.078107), (125,-0.087193), (126,0.185054), (127,0.040655), (128,-0.090738), (129,-0.221205), (130,0.353894), (131,0.211818), (132,0.164958), (133,0.033101), (134,0.397782), (135,0.254310), (136,0.112698), (137,-0.069790), (138,0.309756), (139,0.173717), (140,0.096205), (141,-0.070028), (142,0.185037), (143,0.044814), (144,-0.025265), (145,-0.157591), (146,0.380351), (147,0.215514), (148,0.182592), (149,0.017749), (150,0.385686), (151,0.223173), (152,-0.010874), (153,-0.084210), (154,0.163886), (155,0.180199), (156,0.073427), (157,0.043754), (158,-0.152209), (159,0.118647), (160,-0.040617), (161,-0.100013), (162,0.109529), (163,0.287951), (164,0.134260), (165,0.069754), (166,-0.000325), (167,0.264489), (168,0.046703), (169,-0.043820), (170,0.218214), (171,0.228491), (172,0.073867), (173,0.041877), (174,-0.146654), (175,0.111661), (176,-0.028092), (177,-0.065660), (178,0.181045), (179,0.305585), (180,0.156071), (181,0.084132), (182,-0.006385), (183,0.286300), (184,-0.015098), (185,-0.071708), (186,0.207508), (187,0.191310), (188,0.027864), (189,-0.036642), (190,-0.187084), (191,0.105138), (192,-0.075954), (193,-0.146040), (194,0.113208), (195,0.254936), (196,0.105421), (197,0.038592), (198,-0.032883), (199,0.243546), (200,0.022968), (201,0.004911), (202,0.261372), (203,0.303233), (204,0.137927), (205,0.123119), (206,-0.069125), (207,0.193372), (208,0.057796), (209,0.009082), (210,0.212588), (211,0.352920), (212,0.186224), (213,0.131473), (214,0.129672), (215,0.379627), (216,-0.043936), (217,-0.088937), (218,0.151725), (219,0.132278), (220,-0.002371), (221,-0.068273), (222,-0.195954), (223,0.081872), (224,-0.089934), (225,-0.140508), (226,0.082973), (227,0.213086), (228,0.039890), (229,0.040411), (230,-0.052435), (231,0.265340), (232,0.096784), (233,0.033204), (234,0.267831), (235,0.291577), (236,0.095156), (237,0.061764), (238,-0.126297), (239,0.156175), (240,0.012233), (241,-0.023939), (242,0.229736), (243,0.375177), (244,0.186183), (245,0.141188), (246,0.080859), (247,0.357751), (248,0.186878), (249,0.133518), (250,0.373254), (251,0.376099), (252,0.202433), (253,0.158358), (254,-0.036672), (255,0.268561), (256,0.087926), (257,0.030852), (258,0.278948), (259,0.440188), (260,0.286033), (261,0.208052), (262,0.142613), (263,0.429731), (264,0.084201), (265,0.025731), (266,0.264540), (267,0.290609), (268,0.134595), (269,0.092381), (270,-0.114722), (271,0.171926), (272,0.006156), (273,-0.030943), (274,0.206001), (275,0.371423), (276,0.183819), (277,0.145324), (278,0.075245), (279,0.351211), (280,0.258365), (281,0.093528), (282,0.119133), (283,0.334249), (284,0.292040), (285,0.124411), (286,0.391554), (287,0.213242), (288,0.164065), (289,0.000154), (290,0.187869), (291,0.429928), (292,0.372848), (293,0.199652), (294,0.508598), (295,0.413429), (296,0.091593), (297,-0.051879), (298,0.365294), (299,0.217176), (300,0.143377), (301,-0.005668), (302,0.256366), (303,0.108248), (304,0.052565), (305,-0.098804), (306,0.418237), (307,0.278948), (308,0.235337), (309,0.060281), (310,0.411030), (311,0.243407), (312,0.105044), (313,-0.049573), (314,0.329510), (315,0.212049), (316,0.153579), (317,-0.000112), (318,0.287469), (319,0.119376), (320,0.065553), (321,-0.108576), (322,0.425183), (323,0.327696), (324,0.241819), (325,0.076982), (326,0.472791), (327,0.326532), (328,0.157512), (329,0.020540), (330,0.427494), (331,0.279846), (332,0.199078), (333,0.037027), (334,0.280477), (335,0.122146), (336,0.058566), (337,-0.085375), (338,0.447457), (339,0.311418), (340,0.252484), (341,0.105763), (342,0.479273), (343,0.323259), (344,0.334926), (345,0.143151), (346,0.138563), (347,0.430321), (348,0.351877), (349,0.192149), (350,0.449537), (351,0.274475), (352,0.222511), (353,0.041876), (354,0.238419), (355,0.460967), (356,0.400174), (357,0.258098), (358,0.517339), (359,0.444937), (360,0.185806), (361,0.023755), (362,0.426527), (363,0.283055), (364,0.235267), (365,0.096441), (366,0.332927), (367,0.186206), (368,0.120303), (369,-0.011096), (370,0.507341), (371,0.338784), (372,0.282637), (373,0.159603), (374,0.509426), (375,0.329254), (376,0.116572), (377,-0.013425), (378,0.384237), (379,0.253770), (380,0.196697), (381,0.034177), (382,0.305503), (383,0.109076), (384,0.003230), (385,-0.022259), (386,0.191929), (387,0.329938), (388,0.150236), (389,0.086193), (390,0.031906), (391,0.333883), (392,0.078002), (393,0.051585), (394,0.253695), (395,0.279301), (396,0.145578), (397,0.076426), (398,-0.106526), (399,0.180122), (400,0.034791), (401,-0.038075), (402,0.197478), (403,0.357785), (404,0.204094), (405,0.127509), (406,0.068113), (407,0.364053), (408,-0.006554), (409,-0.007429), (410,0.209545), (411,0.230968), (412,0.091216), (413,0.037392), (414,-0.151139), (415,0.146198), (416,-0.033041), (417,-0.092443), (418,0.174700), (419,0.296454), (420,0.109319), (421,0.059678), (422,0.022110), (423,0.319904), (424,0.214058), (425,0.058971), (426,0.375350), (427,0.197507), (428,0.218004), (429,0.073598), (430,0.023494), (431,-0.131130), (432,0.159701), (433,0.032954), (434,0.360016), (435,0.203532), (436,0.330401), (437,0.185070), (438,0.187451), (439,0.039332), (440,0.150867), (441,-0.023726), (442,0.299153), (443,0.138962), (444,0.146910), (445,-0.020713), (446,-0.101481), (447,-0.248203), (448,0.013368), (449,-0.116172), (450,0.214139), (451,0.090178), (452,0.218901), (453,0.136744), (454,0.160489), (455,0.003542), (456,0.283228), (457,0.112348), (458,0.473317), (459,0.309876), (460,0.319684), (461,0.160883), (462,0.075475), (463,-0.089831), (464,0.175453), (465,0.013402), (466,0.359505), (467,0.201174), (468,0.347543), (469,0.200357), (470,0.223170), (471,0.054620), (472,0.053282), (473,-0.105055), (474,0.252663), (475,0.105008), (476,0.125504), (477,-0.037473), (478,-0.076901), (479,-0.252890), (480,0.012394), (481,-0.173808), (482,0.189947), (483,0.026500), (484,0.176588), (485,0.035439), (486,0.060581), (487,-0.086141), (488,0.220483), (489,0.045884), (490,0.409175), (491,0.250381), (492,0.230928), (493,0.058188), (494,-0.007244), (495,-0.140034), (496,0.129426), (497,-0.054452), (498,0.301406), (499,0.156075), (500,0.294090), (501,0.160837), (502,0.193405), (503,0.025782), (504,0.384427), (505,0.228876), (506,0.185735), (507,0.419898), (508,0.460363), (509,0.311318), (510,0.276542), (511,0.081512), (512,0.337966), (513,0.194958), (514,0.134635), (515,0.368328), (516,0.535604), (517,0.367981), (518,0.338772), (519,0.284485), (520,0.376508), (521,0.213061), (522,0.128580), (523,0.398973), (524,0.418079), (525,0.262065), (526,0.238892), (527,0.031326), (528,0.295677), (529,0.138272), (530,0.103954), (531,0.342763), (532,0.482632), (533,0.301533), (534,0.257465), (535,0.195746), (536,0.255258), (537,0.223263), (538,0.081187), (539,0.461661), (540,0.318188), (541,0.255542), (542,0.119503), (543,0.389890), (544,0.255710), (545,0.179588), (546,0.021251), (547,0.549444), (548,0.391106), (549,0.338673), (550,0.154794), (551,0.558029), (552,0.147471), (553,0.086215), (554,0.316665), (555,0.314863), (556,0.180677), (557,0.085514), (558,-0.093725), (559,0.178992), (560,0.015082), (561,-0.047571), (562,0.208427), (563,0.392421), (564,0.223865), (565,0.144957), (566,0.112035), (567,0.374995), (568,0.235243), (569,0.187455), (570,0.048629), (571,0.440718), (572,0.273095), (573,0.231344), (574,0.075799), (575,0.350832), (576,0.211080), (577,0.137745), (578,-0.011764), (579,0.521996), (580,0.346476), (581,0.314944), (582,0.189587), (583,0.559384), (584,0.307216), (585,0.227845), (586,0.062081), (587,0.478785), (588,0.305588), (589,0.279166), (590,0.121761), (591,0.354528), (592,0.225921), (593,0.175811), (594,0.019797), (595,0.547520), (596,0.393829), (597,0.309817), (598,0.163559), (599,0.518485), (600,0.270036), (601,0.221785), (602,0.062521), (603,0.481554), (604,0.320893), (605,0.251741), (606,0.098513), (607,0.361480), (608,0.219398), (609,0.132594), (610,-0.001585), (611,0.534497), (612,0.378019), (613,0.324659), (614,0.174681), (615,0.557021), (616,0.211954), (617,0.130729), (618,0.391367), (619,0.372377), (620,0.192675), (621,0.176941), (622,-0.016700), (623,0.255090), (624,0.061913), (625,0.036886), (626,0.301707), (627,0.457367), (628,0.311578), (629,0.237310), (630,0.200212), (631,0.489646), (632,0.146909), (633,0.111201), (634,0.349077), (635,0.386292), (636,0.223308), (637,0.181563), (638,-0.011144), (639,0.277364), (640,-0.156418), (641,-0.243685), (642,-0.017888), (643,0.138243), (644,-0.006156), (645,-0.044188), (646,-0.090122), (647,0.198856), (648,-0.107194), (649,-0.160555), (650,0.062000), (651,0.096891), (652,-0.086524), (653,-0.151036), (654,-0.322842), (655,-0.045017), (656,-0.213573), (657,-0.220484), (658,0.014612), (659,0.159127), (660,0.017508), (661,-0.053967), (662,-0.135662), (663,0.144024), (664,0.157551), (665,-0.010079), (666,-0.063902), (667,0.145646), (668,0.159636), (669,0.001763), (670,-0.002826), (671,-0.201569), (672,0.072074), (673,-0.064429), (674,-0.117790), (675,0.135415), (676,0.278534), (677,0.124843), (678,0.069159), (679,-0.011602), (680,0.123157), (681,-0.037503), (682,0.320215), (683,0.148872), (684,0.156363), (685,-0.009407), (686,-0.084595), (687,-0.222031), (688,0.058581), (689,-0.088604), (690,0.267718), (691,0.108454), (692,0.209306), (693,0.055615), (694,0.103976), (695,-0.065971), (696,-0.054767), (697,-0.213098), (698,0.146937), (699,-0.016503), (700,0.032791), (701,-0.124157), (702,-0.241618), (703,-0.379511), (704,-0.119806), (705,-0.267455), (706,0.058210), (707,-0.102450), (708,0.037425), (709,-0.091652), (710,-0.049327), (711,-0.221597), (712,0.040437), (713,-0.123936), (714,0.201729), (715,0.048501), (716,0.088972), (717,-0.068439), (718,-0.147810), (719,-0.294995), (720,-0.007414), (721,-0.148569), (722,0.177102), (723,0.008546), (724,0.145165), (725,0.013772), (726,0.070961), (727,-0.118960), (728,0.109161), (729,-0.011087), (730,-0.060264), (731,0.171576), (732,0.186956), (733,0.027692), (734,-0.033564), (735,-0.185859), (736,0.092893), (737,-0.084486), (738,-0.170363), (739,0.094458), (740,0.257087), (741,0.069953), (742,-0.004772), (743,-0.055346), (744,0.177884), (745,0.042308), (746,0.039116), (747,0.256091), (748,0.324426), (749,0.158199), (750,0.090900), (751,-0.079046), (752,0.209462), (753,0.040906), (754,-0.017100), (755,0.206844), (756,0.366224), (757,0.237617), (758,0.176824), (759,0.083514), (760,0.352054), (761,0.186284), (762,0.115272), (763,0.393561), (764,0.397802), (765,0.210198), (766,0.129900), (767,-0.049802), (768,0.241029), (769,0.109166), (770,0.070208), (771,0.308084), (772,0.450276), (773,0.284042), (774,0.225573), (775,0.145275), (776,0.275851), (777,0.102655), (778,0.065550), (779,0.304359), (780,0.334141), (781,0.143757), (782,0.100152), (783,-0.053539), (784,0.231250), (785,0.056657), (786,-0.010172), (787,0.220741), (788,0.388011), (789,0.253831), (790,0.193502), (791,0.129929), (792,0.184325), (793,0.130038), (794,-0.042231), (795,0.380515), (796,0.227287), (797,0.163245), (798,0.016059), (799,0.256259), (800,0.091885), (801,0.026909), (802,-0.104020), (803,0.442751), (804,0.265365), (805,0.211542), (806,0.075039), (807,0.428574), (808,0.145755), (809,0.110047), (810,-0.032035), (811,0.354480), (812,0.211008), (813,0.147435), (814,-0.021121), (815,0.227438), (816,0.068174), (817,0.021783), (818,-0.099398), (819,0.438544), (820,0.228185), (821,0.205482), (822,0.071765), (823,0.435990), (824,0.182895), (825,0.095627), (826,-0.058527), (827,0.372115), (828,0.228179), (829,0.165990), (830,-0.011389), (831,0.259931), (832,0.096491), (833,0.031052), (834,-0.091056), (835,0.426448), (836,0.294592), (837,0.224970), (838,0.105192), (839,0.433180), (840,0.145714), (841,0.104896), (842,-0.078989), (843,0.363732), (844,0.235589), (845,0.186411), (846,0.017855), (847,0.292894), (848,0.093217), (849,0.065405), (850,-0.081787), (851,0.473343), (852,0.323835), (853,0.244464), (854,0.104705), (855,0.496794), (856,0.214438), (857,0.148072), (858,-0.003759), (859,0.343277), (860,0.249040), (861,0.183138), (862,0.020624), (863,0.267323), (864,0.123851), (865,0.061668), (866,-0.060439), (867,0.489581), (868,0.316842), (869,0.234685), (870,0.067061), (871,0.451254), (872,0.116876), (873,0.073272), (874,0.302789), (875,0.313529), (876,0.164014), (877,0.112977), (878,-0.046750), (879,0.224106), (880,0.078775), (881,0.027274), (882,0.268870), (883,0.410598), (884,0.222994), (885,0.149665), (886,0.090262), (887,0.362052), (888,-0.052688), (889,-0.101403), (890,0.176423), (891,0.176481), (892,0.024650), (893,-0.040326), (894,-0.227924), (895,0.039683), (896,-0.028543), (897,-0.083293), (898,-0.230021), (899,0.316750), (900,0.174668), (901,0.128740), (902,-0.020768), (903,0.308147), (904,0.089428), (905,0.006344), (906,-0.117623), (907,0.285618), (908,0.139822), (909,0.056732), (910,-0.092777), (911,0.153929), (912,-0.010445), (913,-0.041977), (914,-0.184053), (915,0.378504), (916,0.188119), (917,0.144515), (918,-0.042157), (919,0.339713), (920,0.201351), (921,0.040227), (922,-0.026602), (923,0.247041), (924,0.273573), (925,0.087372), (926,0.036334), (927,-0.151733), (928,0.102405), (929,-0.038744), (930,-0.120439), (931,0.143449), (932,0.288427), (933,0.123126), (934,0.082308), (935,-0.000313), (936,-0.010010), (937,-0.137691), (938,0.186584), (939,0.058904), (940,0.074284), (941,-0.079870), (942,-0.170850), (943,-0.325474), (944,-0.075050), (945,-0.191121), (946,0.151269), (947,-0.017287), (948,0.131874), (949,-0.026463), (950,0.012611), (951,-0.139684), (952,0.114454), (953,-0.048529), (954,-0.156698), (955,0.103007), (956,0.114680), (957,-0.041797), (958,-0.117456), (959,-0.272073), (960,0.018288), (961,-0.141439), (962,-0.210591), (963,0.032395), (964,0.175050), (965,0.054339), (966,0.003765), (967,-0.072350), (968,0.197573), (969,0.048528), (970,0.027222), (971,0.264635), (972,0.267009), (973,0.104959), (974,0.036270), (975,-0.158297), (976,0.112566), (977,-0.022547), (978,-0.050823), (979,0.139671), (980,0.297661), (981,0.112849), (982,0.065989), (983,-0.010596), (984,0.132059), (985,-0.033705), (986,-0.052695), (987,0.183328), (988,0.164802), (989,0.029226), (990,-0.020415), (991,-0.195941), (992,0.088391), (993,-0.093634), (994,-0.153964), (995,0.078340), (996,0.214958), (997,0.058944), (998,0.006980), (999,-0.031985), (1000,0.240732), (1001,0.063816), (1002,0.003023), (1003,0.247405), (1004,0.274401), (1005,0.126753), (1006,0.064100), (1007,-0.117462), (1008,0.129707), (1009,-0.028161), (1010,-0.066662), (1011,0.160538), (1012,0.340350), (1013,0.177836), (1014,0.150487), (1015,0.077615), (1016,0.250934), (1017,0.089347), (1018,0.036913), (1019,0.283618), (1020,0.279957), (1021,0.138345), (1022,0.057577), (1023,-0.146740), (1024,0.131080), (1025,-0.012856), (1026,-0.075039), (1027,0.164234), (1028,0.288774), (1029,0.152735), (1030,0.097051), (1031,0.054837), (1032,0.206321), (1033,0.060526), (1034,-0.001194), (1035,0.239469), (1036,0.256715), (1037,0.108134), (1038,0.037585), (1039,-0.165342), (1040,0.106905), (1041,-0.034244), (1042,-0.077849), (1043,0.116835), (1044,0.242301), (1045,0.092330), (1046,0.039896), (1047,-0.001849), (1048,0.081352), (1049,0.023809), (1050,-0.129419), (1051,0.272895), (1052,0.131746), (1053,0.027291), (1054,-0.072055), (1055,0.164894), (1056,0.012593), (1057,-0.063528), (1058,-0.200031), (1059,0.331411), (1060,0.189793), (1061,0.135969), (1062,0.001789), (1063,0.350215), (1064,0.144502), (1065,0.121336), (1066,-0.043507), (1067,0.343478), (1068,0.155410), (1069,0.098800), (1070,-0.063713), (1071,0.190418), (1072,0.059025), (1073,-0.003164), (1074,-0.157782), (1075,0.380623), (1076,0.284070), (1077,0.241392), (1078,0.096060), (1079,0.428694), (1080,0.096640), (1081,0.032127), (1082,-0.129923), (1083,0.246374), (1084,0.102902), (1085,0.065803), (1086,-0.092998), (1087,0.131410), (1088,-0.036220), (1089,-0.083538), (1090,-0.229333), (1091,0.326724), (1092,0.144699), (1093,0.074614), (1094,-0.102765), (1095,0.255880), (1096,0.009760), (1097,-0.011553), (1098,-0.149452), (1099,0.296519), (1100,0.141901), (1101,0.066712), (1102,-0.068864), (1103,0.173195), (1104,0.070593), (1105,0.015843), (1106,-0.146207), (1107,0.411703), (1108,0.267768), (1109,0.181897), (1110,-0.013604), (1111,0.358053), (1112,0.121213), (1113,0.026983), (1114,-0.136464), (1115,0.277923), (1116,0.137237), (1117,0.029062), (1118,-0.104654), (1119,0.147161), (1120,0.010658), (1121,-0.051531), (1122,-0.193607), (1123,0.329007), (1124,0.177639), (1125,0.116846), (1126,0.014250), (1127,0.384041), (1128,0.006927), (1129,-0.047823), (1130,0.191913), (1131,0.222158), (1132,0.050822), (1133,0.005357), (1134,-0.176204), (1135,0.082573), (1136,-0.084123), (1137,-0.125868), (1138,0.114331), (1139,0.267205), (1140,0.113978), (1141,0.053654), (1142,-0.030826), (1143,0.251176), (1144,0.093772), (1145,0.025546), (1146,-0.094701), (1147,0.310393), (1148,0.146952), (1149,0.107524), (1150,-0.041521), (1151,0.216794), (1152,-0.080427), (1153,-0.144007), (1154,-0.312557), (1155,0.236068), (1156,0.053579), (1157,0.017864), (1158,-0.117242), (1159,0.237683), (1160,0.079816), (1161,-0.134263), (1162,-0.182977), (1163,0.065588), (1164,0.072609), (1165,-0.076899), (1166,-0.137229), (1167,-0.331333), (1168,-0.066049), (1169,-0.198369), (1170,-0.227115), (1171,0.042815), (1172,0.173861), (1173,0.024346), (1174,-0.023904), (1175,-0.099093), (1176,-0.030288), (1177,-0.179802), (1178,-0.248491), (1179,-0.007359), (1180,0.005241), (1181,-0.176784), (1182,-0.238510), (1183,-0.424248), (1184,-0.150605), (1185,-0.305686), (1186,-0.367876), (1187,-0.134176), (1188,0.022881), (1189,-0.116414), (1190,-0.145154), (1191,-0.189691), (1192,-0.063292), (1193,-0.209550), (1194,0.113328), (1195,-0.068690), (1196,-0.054700), (1197,-0.194922), (1198,-0.272434), (1199,-0.414979), (1200,-0.151092), (1201,-0.298277), (1202,0.047363), (1203,-0.089604), (1204,0.040046), (1205,-0.147552), (1206,-0.149817), (1207,-0.303045), (1208,-0.023366), (1209,-0.184489), (1210,-0.247136), (1211,-0.000900), (1212,0.004267), (1213,-0.128522), (1214,-0.197211), (1215,-0.316989), (1216,-0.026164), (1217,-0.211439), (1218,-0.261543), (1219,-0.020880), (1220,0.124098), (1221,-0.048172), (1222,-0.077381), (1223,-0.148856), (1224,0.094600), (1225,-0.072567), (1226,-0.118494), (1227,0.069220), (1228,0.060918), (1229,-0.075121), (1230,-0.127091), (1231,-0.293325), (1232,-0.016425), (1233,-0.169653), (1234,-0.191430), (1235,0.042270), (1236,0.206296), (1237,0.125529), (1238,0.055443), (1239,-0.026251), (1240,0.006324), (1241,-0.162696), (1242,-0.252286), (1243,0.029716), (1244,0.026525), (1245,-0.097442), (1246,-0.164735), (1247,-0.356516), (1248,-0.067544), (1249,-0.262105), (1250,-0.337300), (1251,-0.101277), (1252,0.041841), (1253,-0.134148), (1254,-0.138266), (1255,-0.255727), (1256,0.051823), (1257,-0.129739), (1258,-0.151509), (1259,0.118414), (1260,0.135661), (1261,-0.033359), (1262,-0.058385), (1263,-0.252026), (1264,0.024873), (1265,-0.165981), (1266,-0.217018), (1267,0.030151), (1268,0.202536), (1269,0.029340), (1270,-0.004515), (1271,-0.100605), (1272,0.140058), (1273,-0.035931), (1274,-0.104620), (1275,0.129543), (1276,0.148643), (1277,-0.006438), (1278,-0.035647), (1279,-0.220922), (1280,0.026246), (1281,-0.138127), (1282,-0.177092), (1283,0.086338), (1284,0.230383), (1285,0.076692), (1286,-0.007319), (1287,-0.071368), (1288,0.094981), (1289,-0.056387), (1290,-0.119039), (1291,0.139745), (1292,0.150949), (1293,-0.039436), (1294,-0.058889), (1295,-0.264602), (1296,-0.027653), (1297,-0.173448), (1298,-0.239350), (1299,-0.001937), (1300,0.139791), (1301,0.004215), (1302,-0.039859), (1303,-0.110865), (1304,0.120505), (1305,0.086657), (1306,-0.079113), (1307,-0.052581), (1308,0.197374), (1309,0.142160), (1310,-0.020823), (1311,0.261186), (1312,0.051290), (1313,0.014185), (1314,-0.161804), (1315,-0.026112), (1316,0.190863), (1317,0.122174), (1318,-0.031517), (1319,0.230053), (1320,-0.075527), (1321,-0.136783), (1322,-0.289548), (1323,0.095578), (1324,-0.026066), (1325,-0.106834), (1326,-0.215002), (1327,0.045635), (1328,-0.076002), (1329,-0.128436), (1330,-0.285840), (1331,0.259534), (1332,0.089118), (1333,0.005101), (1334,-0.172278), (1335,0.192410), (1336,-0.090416), (1337,-0.118692), (1338,-0.271920), (1339,0.159192), (1340,-0.007505), (1341,-0.065975), (1342,-0.208520), (1343,0.023784), (1344,-0.108536), (1345,-0.134496), (1346,-0.306765), (1347,0.240933), (1348,0.108606), (1349,0.078007), (1350,-0.104018), (1351,0.239299), (1352,0.047524), (1353,-0.014665), (1354,-0.145595), (1355,0.228379), (1356,0.036598), (1357,-0.024659), (1358,-0.199251), (1359,0.023303), (1360,-0.137357), (1361,-0.162847), (1362,-0.313288), (1363,0.224654), (1364,0.132277), (1365,0.076130), (1366,-0.093353), (1367,0.262043), (1368,0.121820), (1369,0.072643), (1370,-0.067116), (1371,-0.056839), (1372,0.168495), (1373,0.129073), (1374,-0.018118), (1375,0.241593), (1376,0.044702), (1377,-0.017481), (1378,-0.185574), (1379,-0.046168), (1380,0.206110), (1381,0.184803), (1382,0.014850), (1383,0.278744), (1384,0.002888), (1385,-0.154517), (1386,0.224567), (1387,0.074589), (1388,0.074647), (1389,-0.099013), (1390,-0.194646), (1391,-0.341368), (1392,-0.037994), (1393,-0.213983), (1394,0.084281), (1395,-0.064301), (1396,0.093220), (1397,-0.031211), (1398,-0.042768), (1399,-0.196453), (1400,-0.042652), (1401,-0.084867), (1402,-0.251093), (1403,0.188371), (1404,0.061161), (1405,-0.001492), (1406,-0.137068), (1407,0.080840), (1408,-0.037554), (1409,-0.204251), (1410,-0.248782), (1411,-0.003010), (1412,0.141505), (1413,-0.033551), (1414,-0.079015), (1415,-0.163033), (1416,-0.044066), (1417,-0.194507), (1418,-0.239971), (1419,0.006271), (1420,0.030943), (1421,-0.126924), (1422,-0.185857), (1423,-0.362773), (1424,-0.057546), (1425,-0.226566), (1426,-0.251129), (1427,-0.024398), (1428,0.107574), (1429,-0.031251), (1430,-0.077179), (1431,-0.150978), (1432,0.027914), (1433,-0.120204), (1434,-0.151737), (1435,0.094042), (1436,0.093167), (1437,-0.082352), (1438,-0.125963), (1439,-0.316811), (1440,-0.058033), (1441,-0.189426), (1442,-0.227921), (1443,0.031326), (1444,0.180944), (1445,0.027723), (1446,-0.043289), (1447,-0.103619), (1448,-0.406413), (1449,-0.134623), (1450,0.109752), (1451,0.050819), (1452,-0.095903), (1453,-0.081449), (1454,-0.281589), (1455,-0.368856), (1456,-0.542053), (1457,-0.265623), (1458,-0.057008), (1459,-0.067632), (1460,-0.212964), (1461,-0.053584), (1462,-0.119950), (1463,-0.174706), (1464,-0.327471), (1465,-0.028274), (1466,-0.200549), (1467,0.107007), (1468,-0.033679), (1469,-0.002500), (1470,-0.152478), (1471,-0.227203), (1472,-0.354883), (1473,-0.092850), (1474,-0.275808), (1475,0.093526), (1476,-0.096395), (1477,0.052296), (1478,-0.089316), (1479,-0.058137), (1480,-0.237376), (1481,0.033017), (1482,-0.164337), (1483,0.208710), (1484,0.074994), (1485,0.122428), (1486,-0.056347), (1487,-0.139902), (1488,-0.277331), (1489,0.004671), (1490,-0.154129), (1491,0.189187), (1492,0.009022), (1493,0.184194), (1494,0.048154), (1495,0.070974), (1496,-0.281989), (1497,-0.018565), (1498,-0.195011), (1499,0.175243), (1500,0.018302), (1501,0.053664), (1502,-0.120002), (1503,-0.206343), (1504,-0.322871), (1505,-0.044581), (1506,-0.187590), (1507,0.121356), (1508,-0.015153), (1509,0.091742), (1510,-0.047554), (1511,-0.013589), (1512,-0.175176), (1513,0.126338), (1514,-0.023634), (1515,0.298781), (1516,0.109324), (1517,0.126100), (1518,-0.032700), (1519,-0.115321), (1520,-0.268549), (1521,0.006027), (1522,-0.128622), (1523,0.243498), (1524,0.084228), (1525,0.247327), (1526,0.078771), (1527,0.147569), (1528,-0.137103), (1529,0.127247), (1530,-0.042699), (1531,0.302014), (1532,0.134384), (1533,0.157204), (1534,0.015591), (1535,-0.108376), (1536,-0.235123), (1537,0.035270), (1538,-0.107738), (1539,0.264839), (1540,0.113008), (1541,0.274711), (1542,0.072248), (1543,0.115035), (1544,-0.195191), (1545,0.067776), (1546,-0.125865), (1547,0.245786), (1548,0.114392), (1549,0.106091), (1550,-0.059679), (1551,-0.182713), (1552,-0.308070), (1553,-0.015385), (1554,-0.165357), (1555,0.160308), (1556,0.008014), (1557,0.150669), (1558,0.028561), (1559,0.061136), (1560,0.281361), (1561,0.146255), (1562,0.079419), (1563,-0.059407), (1564,0.301098), (1565,0.140908), (1566,0.070822), (1567,-0.075436), (1568,0.196817), (1569,0.009682), (1570,-0.053434), (1571,-0.221990), (1572,0.328494), (1573,0.169230), (1574,0.152100), (1575,-0.003451), (1576,0.209810), (1577,0.053796), (1578,-0.015819), (1579,0.252714), (1580,0.242090), (1581,0.080033), (1582,-0.002125), (1583,-0.153956), (1584,0.108541), (1585,-0.047473), (1586,-0.092937), (1587,0.138903), (1588,0.271339), (1589,0.123227), (1590,0.095878), (1591,0.000245), (1592,0.114102), (1593,-0.041912), (1594,-0.099449), (1595,0.180700), (1596,0.227671), (1597,0.065614), (1598,-0.018867), (1599,-0.228293), (1600,0.061605), (1601,-0.100909), (1602,-0.137087), (1603,0.078035), (1604,0.235555), (1605,0.079077), (1606,-0.030024), (1607,-0.095927), (1608,0.098293), (1609,-0.025210), (1610,-0.080888), (1611,0.158849), (1612,0.156114), (1613,0.034013), (1614,-0.013775), (1615,-0.212988), (1616,0.065301), (1617,-0.124157), (1618,-0.154292), (1619,0.071048), (1620,0.257829), (1621,0.086950), (1622,0.045668), (1623,-0.038813), (1624,0.259915), (1625,0.092291), (1626,0.052863), (1627,-0.087822), (1628,0.321455), (1629,0.188202), (1630,0.119513), (1631,-0.021173), (1632,0.245507), (1633,0.078811), (1634,0.049138), (1635,-0.108736), (1636,0.422243), (1637,0.269016), (1638,0.214259), (1639,0.049422), (1640,0.036938), (1641,-0.082846), (1642,0.237246), (1643,0.090524), (1644,0.087332), (1645,-0.084943), (1646,-0.182430), (1647,-0.351449), (1648,-0.066654), (1649,-0.201767), (1650,0.179176), (1651,0.025022), (1652,0.169536), (1653,0.036283), (1654,0.065602), (1655,-0.089485), (1656,0.154897), (1657,-0.005757), (1658,-0.054478), (1659,0.192691), (1660,0.227119), (1661,-0.009714), (1662,-0.054715), (1663,-0.217229), (1664,-0.105694), (1665,-0.256129), (1666,-0.316459), (1667,-0.086478), (1668,0.076151), (1669,-0.069644), (1670,-0.135546), (1671,-0.189833), (1672,-0.008162), (1673,-0.193900), (1674,-0.247260), (1675,0.013377), (1676,0.045952), (1677,-0.117495), (1678,-0.205695), (1679,-0.323619), (1680,-0.090383), (1681,-0.259403), (1682,-0.327628), (1683,-0.080459), (1684,0.080774), (1685,-0.090562), (1686,-0.135563), (1687,-0.208435), (1688,-0.450378), (1689,-0.157687), (1690,-0.284904), (1691,0.073741), (1692,-0.114784), (1693,-0.130987), (1694,-0.267490), (1695,-0.334789), (1696,-0.482901), (1697,-0.191606), (1698,-0.353663), (1699,-0.018705), (1700,-0.242533), (1701,-0.087800), (1702,-0.229412), (1703,-0.179655), (1704,-0.368186), (1705,-0.090360), (1706,-0.256593), (1707,0.116917), (1708,-0.029805), (1709,-0.000016), (1710,-0.189944), (1711,-0.272565), (1712,-0.431829), (1713,-0.153540), (1714,-0.286793), (1715,0.046305), (1716,-0.120855), (1717,0.014367), (1718,-0.174157), (1719,-0.123937), (1720,-0.442060), (1721,-0.157265), (1722,-0.310492), (1723,0.042580), (1724,-0.093459), (1725,-0.072963), (1726,-0.222008), (1727,-0.365480), (1728,-0.446248), (1729,-0.181897), (1730,-0.356490), (1731,-0.010844), (1732,-0.121805), (1733,0.041758), (1734,-0.107294), (1735,-0.086334), (1736,-0.303193), (1737,-0.054634), (1738,-0.188814), (1739,0.160539), (1740,0.030542), (1741,-0.012599), (1742,-0.181619), (1743,-0.226157), (1744,-0.403536), (1745,-0.123387), (1746,-0.258499), (1747,0.058806), (1748,-0.101384), (1749,0.069605), (1750,-0.074794), (1751,-0.025970), (1752,-0.452320), (1753,-0.209327), (1754,-0.359769), (1755,-0.014129), (1756,-0.143669), (1757,-0.137568), (1758,-0.256426), (1759,-0.342766), (1760,-0.500634), (1761,-0.217698), (1762,-0.368140), (1763,0.001651), (1764,-0.169685), (1765,-0.052578), (1766,-0.209519), (1767,-0.175554), (1768,-0.332501), (1769,-0.091368), (1770,-0.239487), (1771,0.085715), (1772,-0.096310), (1773,-0.074418), (1774,-0.180733), (1775,-0.245702), (1776,-0.394284), (1777,-0.132720), (1778,-0.272472), (1779,0.070844), (1780,-0.068915), (1781,0.101611), (1782,-0.081804), (1783,-0.060381), (1784,-0.216859), (1785,0.084655), (1786,-0.103406), (1787,0.214363), (1788,0.081573), (1789,0.078381), (1790,-0.127338), (1791,-0.229934), (1792,-0.321848), (1793,-0.046345), (1794,-0.201426), (1795,0.125635), (1796,-0.023879), (1797,0.139220), (1798,-0.021903), (1799,0.032500), (1800,-0.265655), (1801,0.015427), (1802,-0.157775), (1803,0.169286), (1804,0.047642), (1805,0.037481), (1806,-0.130142), (1807,-0.241567), (1808,-0.421732), (1809,-0.124401), (1810,-0.279946), (1811,0.033640), (1812,-0.118191), (1813,0.023074), (1814,-0.160811), (1815,-0.078537), (1816,0.135651), (1817,-0.049160), (1818,-0.098807), (1819,-0.232060), (1820,0.170254), (1821,0.056506), (1822,-0.025188), (1823,-0.180739), (1824,0.099873), (1825,-0.047312), (1826,-0.105319), (1827,-0.302209), (1828,0.232946), (1829,0.111309), (1830,0.010103), (1831,-0.117114), (1832,-0.033444), (1833,-0.185275), (1834,-0.229813), (1835,0.015960), (1836,0.034133), (1837,-0.094011), (1838,-0.127396), (1839,-0.317781), (1840,-0.047857), (1841,-0.211761), (1842,-0.279060), (1843,-0.032818), (1844,0.126556), (1845,-0.062432), (1846,-0.131584), (1847,-0.196560), (1848,-0.009773), (1849,-0.181579), (1850,-0.244232), (1851,0.016869), (1852,0.028543), (1853,-0.129331), (1854,-0.176186), (1855,-0.340565), (1856,-0.052984), (1857,-0.207138), (1858,-0.246103), (1859,0.008035), (1860,0.133508), (1861,-0.016007), (1862,-0.068434), (1863,-0.146415), (1864,0.044085), (1865,-0.114715), (1866,-0.167612), (1867,0.057259), (1868,0.038275), (1869,-0.121922), (1870,-0.174813), (1871,-0.329900), (1872,-0.027923), (1873,-0.190900), (1874,-0.224756), (1875,0.034492), (1876,0.186903), (1877,-0.001628), (1878,-0.041514), (1879,-0.106489), (1880,0.214536), (1881,0.061308), (1882,-0.022246), (1883,-0.163858), (1884,0.240309), (1885,0.075936), (1886,0.016070), (1887,-0.178028), (1888,0.096078), (1889,-0.044607), (1890,-0.099827), (1891,-0.275347), (1892,0.276528), (1893,0.136775), (1894,0.107103), (1895,-0.068886), (1896,0.070989), (1897,-0.067844), (1898,-0.109589), (1899,0.121319), (1900,0.144138), (1901,-0.011876), (1902,-0.094498), (1903,-0.273273), (1904,0.030101), (1905,-0.082714), (1906,-0.171378), (1907,-0.005498), (1908,0.130657), (1909,-0.006309), (1910,-0.059206), (1911,-0.139974), (1912,-0.015434), (1913,-0.173301), (1914,-0.200651), (1915,0.076712), (1916,0.070264), (1917,-0.091786), (1918,-0.159085), (1919,-0.323922), (1920,-0.218424), (1921,-0.406955), (1922,-0.452882), (1923,-0.221506), (1924,-0.055626), (1925,-0.213030), (1926,-0.236667), (1927,-0.350871), (1928,-0.087911), (1929,-0.243925), (1930,-0.289389), (1931,-0.034788), (1932,-0.017548), (1933,-0.186568), (1934,-0.234819), (1935,-0.415447), (1936,-0.113007), (1937,-0.223035), (1938,-0.299620), (1939,-0.082645), (1940,0.081844), (1941,-0.070914), (1942,-0.131243), (1943,-0.188323), (1944,-0.439552), (1945,-0.133862), (1946,-0.344685), (1947,-0.028306), (1948,-0.179674), (1949,-0.169397), (1950,-0.291967), (1951,-0.348114), (1952,-0.524103), (1953,-0.268112), (1954,-0.393932), (1955,-0.051079), (1956,-0.174576), (1957,-0.040744), (1958,-0.203727), (1959,-0.208315), (1960,-0.364329), (1961,-0.059560), (1962,-0.251804), (1963,0.094299), (1964,-0.040350), (1965,0.007553), (1966,-0.172612), (1967,-0.259416), (1968,-0.431692), (1969,-0.145037), (1970,-0.291765), (1971,0.080355), (1972,-0.065440), (1973,0.074892), (1974,-0.108060), (1975,-0.063876), (1976,-0.457245), (1977,-0.208223), (1978,-0.365627), (1979,-0.025097), (1980,-0.150917), (1981,-0.150396), (1982,-0.296654), (1983,-0.370453), (1984,-0.548295), (1985,-0.282548), (1986,-0.451568), (1987,-0.079917), (1988,-0.271698), (1989,-0.121140), (1990,-0.275301), (1991,-0.207893), (1992,-0.317451), (1993,-0.005719), (1994,-0.171952), (1995,0.145354), (1996,0.039508), (1997,0.013086), (1998,-0.124350), (1999,-0.214867), (2000,-0.408971), (2001,-0.124640), (2002,-0.281117), (2003,0.075668), (2004,-0.053871), (2005,0.080894), (2006,-0.063974), (2007,-0.045338), (2008,-0.417342), (2009,-0.145089), (2010,-0.318755), (2011,0.006446), (2012,-0.154671), (2013,-0.131395), (2014,-0.312024), (2015,-0.363988), (2016,-0.531617), (2017,-0.248682), (2018,-0.391227), (2019,-0.044191), (2020,-0.183480), (2021,-0.045008), (2022,-0.194980), (2023,-0.156368), (2024,-0.318425), (2025,-0.053605), (2026,-0.211942), (2027,0.122552), (2028,-0.043681), (2029,-0.030618), (2030,-0.187095), (2031,-0.270650), (2032,-0.389964), (2033,-0.136759), (2034,-0.271872), (2035,0.058909), (2036,-0.086423), (2037,0.067848), (2038,-0.084453), (2039,-0.053275), (2040,-0.099666), (2041,0.178160), (2042,-0.001542), (2043,-0.076274), (2044,0.169505), (2045,0.173740), (2046,-0.001316), (2047,-0.048640), (2048,-0.451302), (2049,-0.169757), (2050,0.017951), (2051,-0.022397), (2052,-0.177485), (2053,-0.010672), (2054,-0.073788), (2055,-0.145727), (2056,-0.466636), (2057,-0.188810), (2058,0.037914), (2059,-0.026129), (2060,-0.164954), (2061,-0.166756), (2062,-0.332520), (2063,-0.381240), (2064,-0.526566), (2065,-0.226912), (2066,-0.012260), (2067,-0.039139), (2068,-0.206306), (2069,-0.033457), (2070,-0.112365), (2071,-0.182907), (2072,0.011770), (2073,-0.134952), (2074,-0.206891), (2075,0.027736), (2076,0.025934), (2077,-0.116611), (2078,-0.158819), (2079,-0.325516), (2080,-0.061629), (2081,-0.174444), (2082,-0.221768), (2083,0.004963), (2084,0.163880), (2085,-0.012573), (2086,-0.031563), (2087,-0.114647), (2088,-0.105766), (2089,-0.268750), (2090,0.097798), (2091,-0.073545), (2092,-0.050726), (2093,-0.218819), (2094,-0.336743), (2095,-0.512732), (2096,-0.237229), (2097,-0.395097), (2098,-0.057353), (2099,-0.203148), (2100,-0.038659), (2101,-0.216044), (2102,-0.130984), (2103,-0.267950), (2104,-0.105784), (2105,-0.244616), (2106,0.079659), (2107,-0.065666), (2108,-0.042390), (2109,-0.210477), (2110,-0.305640), (2111,-0.441216), (2112,-0.177792), (2113,-0.333343), (2114,-0.006745), (2115,-0.122810), (2116,-0.004775), (2117,-0.177508), (2118,-0.128215), (2119,-0.308850), (2120,-0.157829), (2121,-0.303161), (2122,0.055484), (2123,-0.117249), (2124,-0.076778), (2125,-0.226756), (2126,-0.297768), (2127,-0.462141), (2128,-0.202894), (2129,-0.333830), (2130,0.010420), (2131,-0.125620), (2132,0.022608), (2133,-0.137119), (2134,-0.111050), (2135,-0.297258), (2136,0.025164), (2137,-0.110413), (2138,-0.173529), (2139,0.060171), (2140,0.076948), (2141,-0.089285), (2142,-0.133823), (2143,-0.312129), (2144,0.007500), (2145,-0.141081), (2146,-0.200948), (2147,0.045294), (2148,0.180517), (2149,0.012893), (2150,-0.031175), (2151,-0.095687), (2152,-0.025022), (2153,-0.192189), (2154,0.125117), (2155,-0.015562), (2156,0.000751), (2157,-0.149690), (2158,-0.223025), (2159,-0.375783), (2160,-0.087745), (2161,-0.237716), (2162,0.114893), (2163,-0.048554), (2164,0.105253), (2165,-0.053084), (2166,-0.017260), (2167,-0.176530), (2168,-0.066849), (2169,-0.229832), (2170,0.126027), (2171,-0.015586), (2172,-0.012278), (2173,-0.144598), (2174,-0.225829), (2175,-0.402281), (2176,-0.421271), (2177,-0.165743), (2178,-0.224213), (2179,-0.365362), (2180,-0.252431), (2181,-0.326693), (2182,-0.391199), (2183,-0.539780), (2184,-0.331165), (2185,-0.101185), (2186,-0.136430), (2187,-0.315205), (2188,-0.323043), (2189,-0.478131), (2190,-0.542173), (2191,-0.703760), (2192,-0.447763), (2193,-0.230324), (2194,-0.285081), (2195,-0.391854), (2196,-0.236656), (2197,-0.306742), (2198,-0.339200), (2199,-0.503574), (2200,-0.660051), (2201,0.035822), (2202,-0.150849), (2203,-0.194454), (2204,-0.345358), (2205,-0.343910), (2206,-0.512930), (2207,-0.535633), (2208,-0.691647), (2209,-0.007389), (2210,-0.169902), (2211,-0.256706), (2212,-0.396929), (2213,-0.156266), (2214,-0.318780), (2215,-0.373536), (2216,-0.555561), (2217,0.148208), (2218,-0.032427), (2219,-0.089500), (2220,-0.279421), (2221,-0.297015), (2222,-0.428878), (2223,-0.511036), (2224,-0.655898), (2225,0.022782), (2226,-0.137872), (2227,-0.204238), (2228,-0.364435), (2229,-0.114017), (2230,-0.250056), (2231,-0.303417), (2232,-0.752527), (2233,-0.055263), (2234,-0.225673), (2235,-0.293898), (2236,-0.446663), (2237,-0.454037), (2238,-0.572425), (2239,-0.647614), (2240,-0.819889), (2241,-0.124948), (2242,-0.294432), (2243,-0.356151), (2244,-0.485691), (2245,-0.261747), (2246,-0.402432), (2247,-0.452073), (2248,-0.651287), (2249,0.043191), (2250,-0.130475), (2251,-0.175006), (2252,-0.329161), (2253,-0.317957), (2254,-0.496269), (2255,-0.568208), (2256,-0.712143), (2257,-0.028818), (2258,-0.195978), (2259,-0.241442), (2260,-0.424394), (2261,-0.128453), (2262,-0.303515), (2263,-0.377777), (2264,-0.686144), (2265,-0.047871), (2266,-0.204349), (2267,-0.233558), (2268,-0.385389), (2269,-0.384868), (2270,-0.549705), (2271,-0.610034), (2272,-0.762329), (2273,-0.060889), (2274,-0.244304), (2275,-0.346436), (2276,-0.515919), (2277,-0.280829), (2278,-0.397827), (2279,-0.469302), (2280,-0.607665), (2281,0.072411), (2282,-0.096139), (2283,-0.173194), (2284,-0.316196), (2285,-0.342155), (2286,-0.496310), (2287,-0.563602), (2288,-0.709398), (2289,-0.046974), (2290,-0.204841), (2291,-0.239623), (2292,-0.417002), (2293,-0.147079), (2294,-0.265003), (2295,-0.316504), (2296,-0.368467), (2297,-0.100397), (2298,0.161630), (2299,0.112453), (2300,-0.019874), (2301,-0.023529), (2302,-0.205090), (2303,-0.288645), (2304,-0.453018), (2305,-0.154291), (2306,0.040393), (2307,-0.038985), (2308,-0.213578), (2309,-0.050015), (2310,-0.105698), (2311,-0.144663), (2312,-0.484150), (2313,-0.208648), (2314,0.040381), (2315,-0.013443), (2316,-0.162494), (2317,-0.174978), (2318,-0.320304), (2319,-0.396889), (2320,-0.549190), (2321,-0.263931), (2322,-0.061358), (2323,-0.078482), (2324,-0.233106), (2325,-0.030990), (2326,-0.088997), (2327,-0.165582), (2328,-0.081454), (2329,-0.232359), (2330,0.078447), (2331,-0.070135), (2332,-0.057534), (2333,-0.219121), (2334,-0.318931), (2335,-0.448471), (2336,-0.198979), (2337,-0.331769), (2338,-0.001921), (2339,-0.133777), (2340,0.013524), (2341,-0.150386), (2342,-0.128500), (2343,-0.272899), (2344,-0.241257), (2345,-0.003844), (2346,-0.050235), (2347,-0.228084), (2348,-0.217343), (2349,-0.397972), (2350,-0.419749), (2351,-0.589232), (2352,-0.265890), (2353,-0.031727), (2354,-0.099946), (2355,-0.294983), (2356,-0.171369), (2357,-0.230766), (2358,-0.324069), (2359,-0.449896), (2360,-0.136767), (2361,-0.241686), (2362,0.054718), (2363,-0.105009), (2364,-0.078477), (2365,-0.239600), (2366,-0.331514), (2367,-0.470803), (2368,-0.181368), (2369,-0.359217), (2370,-0.028436), (2371,-0.203962), (2372,-0.046441), (2373,-0.214528), (2374,-0.144796), (2375,-0.310103), (2376,-0.090341), (2377,-0.219875), (2378,0.105327), (2379,-0.041395), (2380,-0.032051), (2381,-0.199211), (2382,-0.262327), (2383,-0.426237), (2384,-0.118681), (2385,-0.279341), (2386,0.032855), (2387,-0.069278), (2388,0.088706), (2389,-0.067772), (2390,-0.041233), (2391,-0.206539), (2392,-0.055055), (2393,-0.189241), (2394,0.159191), (2395,-0.008902), (2396,0.014381), (2397,-0.148603), (2398,-0.226578), (2399,-0.414176), (2400,-0.130777), (2401,-0.319771), (2402,-0.002466), (2403,-0.129682), (2404,-0.000496), (2405,-0.134213), (2406,-0.120686), (2407,-0.235360), (2408,-0.160519), (2409,0.063425), (2410,0.008205), (2411,-0.161278), (2412,-0.132423), (2413,-0.266602), (2414,-0.333895), (2415,-0.479227), (2416,-0.221376), (2417,0.006282), (2418,0.003090), (2419,-0.183118), (2420,-0.018165), (2421,-0.065489), (2422,-0.137428), (2423,-0.329672), (2424,-0.309639), (2425,-0.054111), (2426,-0.082387), (2427,-0.230969), (2428,-0.209083), (2429,-0.389712), (2430,-0.417524), (2431,-0.608378), (2432,-0.429024), (2433,-0.180002), (2434,-0.217570), (2435,-0.432569), (2436,-0.264830), (2437,-0.353957), (2438,-0.388275), (2439,-0.543356), (2440,-0.377477), (2441,-0.092218), (2442,-0.164627), (2443,-0.326214), (2444,-0.318723), (2445,-0.470091), (2446,-0.558291), (2447,-0.702227), (2448,-0.403036), (2449,-0.168873), (2450,-0.232452), (2451,-0.423764), (2452,-0.293651), (2453,-0.407862), (2454,-0.449143), (2455,-0.586579), (2456,-0.255798), (2457,-0.411349), (2458,-0.086611), (2459,-0.219401), (2460,-0.189149), (2461,-0.339127), (2462,-0.424998), (2463,-0.591231), (2464,-0.314338), (2465,-0.460133), (2466,-0.126103), (2467,-0.307664), (2468,-0.139925), (2469,-0.272245), (2470,-0.231317), (2471,-0.386398), (2472,-0.617659), (2473,0.064740), (2474,-0.092671), (2475,-0.107941), (2476,-0.267669), (2477,-0.274580), (2478,-0.420838), (2479,-0.466766), (2480,-0.638109), (2481,0.001554), (2482,-0.160960), (2483,-0.172517), (2484,-0.343390), (2485,-0.127812), (2486,-0.250382), (2487,-0.319071), (2488,-0.721726), (2489,-0.089033), (2490,-0.238541), (2491,-0.281219), (2492,-0.394497), (2493,-0.428346), (2494,-0.601085), (2495,-0.691602), (2496,-0.848080), (2497,-0.156389), (2498,-0.331914), (2499,-0.373196), (2500,-0.518064), (2501,-0.279255), (2502,-0.410648), (2503,-0.481660), (2504,-0.667405), (2505,-0.016127), (2506,-0.196755), (2507,-0.255225), (2508,-0.406130), (2509,-0.436729), (2510,-0.554190), (2511,-0.640994), (2512,-0.796545), (2513,-0.124365), (2514,-0.293848), (2515,-0.330020), (2516,-0.471633), (2517,-0.210532), (2518,-0.360040), (2519,-0.408754), (2520,-0.584280), (2521,-0.316210), (2522,-0.063931), (2523,-0.128437), (2524,-0.305353), (2525,-0.277431), (2526,-0.467352), (2527,-0.508633), (2528,-0.660465), (2529,-0.405863), (2530,-0.170773), (2531,-0.213451), (2532,-0.378288), (2533,-0.218915), (2534,-0.267629), (2535,-0.334921), (2536,-0.502081), (2537,-0.231225), (2538,0.032199), (2539,-0.004442), (2540,-0.167883), (2541,-0.142747), (2542,-0.335454), (2543,-0.373023), (2544,-0.535073), (2545,-0.238206), (2546,-0.040272), (2547,-0.103388), (2548,-0.262189), (2549,-0.098626), (2550,-0.197972), (2551,-0.242047), (2552,-0.436608), (2553,-0.145783), (2554,0.073522), (2555,0.058715), (2556,-0.126567), (2557,-0.118149), (2558,-0.273231), (2559,-0.365144), (2560,-0.495147), (2561,-0.244265), (2562,-0.008242), (2563,0.018753), (2564,-0.136791), (2565,-0.032226), (2566,-0.101842), (2567,-0.128727), (2568,-0.426412), (2569,-0.139294), (2570,0.073498), (2571,-0.010056), (2572,-0.153528), (2573,-0.135355), (2574,-0.289509), (2575,-0.312213), (2576,-0.487268), (2577,-0.211302), (2578,0.029824), (2579,0.003871), (2580,-0.174905), (2581,-0.019238), (2582,-0.110224), (2583,-0.184949), (2584,-0.106395), (2585,-0.286097), (2586,0.036318), (2587,-0.109014), (2588,-0.091768), (2589,-0.267756), (2590,-0.351304), (2591,-0.499886), (2592,-0.208128), (2593,-0.352063), (2594,-0.018502), (2595,-0.187985), (2596,-0.054153), (2597,-0.190662), (2598,-0.152978), (2599,-0.277408), (2600,-0.138929), (2601,-0.278218), (2602,0.067421), (2603,-0.111818), (2604,-0.093644), (2605,-0.231544), (2606,-0.316488), (2607,-0.444631), (2608,-0.178421), (2609,-0.302851), (2610,0.027930), (2611,-0.141553), (2612,0.011784), (2613,-0.136798), (2614,-0.145105), (2615,-0.313192), (2616,-0.108296), (2617,-0.258267), (2618,0.098055), (2619,-0.065855), (2620,-0.076943), (2621,-0.203233), (2622,-0.329054), (2623,-0.500396), (2624,-0.217461), (2625,-0.378585), (2626,-0.025976), (2627,-0.194995), (2628,-0.037938), (2629,-0.201849), (2630,-0.209686), (2631,-0.335043), (2632,-0.162658), (2633,-0.336324), (2634,-0.036206), (2635,-0.149485), (2636,-0.087649), (2637,-0.273387), (2638,-0.350905), (2639,-0.527357), (2640,-0.248599), (2641,-0.374889), (2642,-0.066406), (2643,-0.190366), (2644,-0.033779), (2645,-0.224627), (2646,-0.184626), (2647,-0.328561), (2648,-0.138524), (2649,-0.296398), (2650,0.065034), (2651,-0.083548), (2652,-0.055156), (2653,-0.224175), (2654,-0.341636), (2655,-0.469310), (2656,-0.210532), (2657,-0.358187), (2658,-0.000005), (2659,-0.177848), (2660,-0.052375), (2661,-0.202816), (2662,-0.183716), (2663,-0.336481), (2664,-0.327130), (2665,-0.078572), (2666,-0.144004), (2667,-0.290263), (2668,-0.276736), (2669,-0.438323), (2670,-0.439661), (2671,-0.625406), (2672,-0.331325), (2673,-0.080437), (2674,-0.135193), (2675,-0.329761), (2676,-0.163875), (2677,-0.182401), (2678,-0.251554), (2679,-0.388520), (2680,-0.384749), (2681,-0.139440), (2682,-0.173289), (2683,-0.343241), (2684,-0.337610), (2685,-0.524745), (2686,-0.556734), (2687,-0.722504), (2688,-0.795839), (2689,-0.126446), (2690,-0.286173), (2691,-0.359508), (2692,-0.506694), (2693,-0.271604), (2694,-0.418789), (2695,-0.514885), (2696,-0.766584), (2697,-0.090221), (2698,-0.205359), (2699,-0.258256), (2700,-0.403125), (2701,-0.454162), (2702,-0.597634), (2703,-0.646812), (2704,-0.804216), (2705,-0.126000), (2706,-0.278295), (2707,-0.328868), (2708,-0.489992), (2709,-0.233537), (2710,-0.365857), (2711,-0.428510), (2712,-0.803301), (2713,-0.138547), (2714,-0.277843), (2715,-0.292187), (2716,-0.429153), (2717,-0.453716), (2718,-0.583719), (2719,-0.652408), (2720,-0.803306), (2721,-0.124164), (2722,-0.263453), (2723,-0.327032), (2724,-0.509057), (2725,-0.277681), (2726,-0.422549), (2727,-0.481946), (2728,-0.402458), (2729,-0.121383), (2730,-0.299231), (2731,-0.354908), (2732,-0.513709), (2733,-0.497865), (2734,-0.633435), (2735,-0.693301), (2736,-0.439163), (2737,-0.174349), (2738,-0.331290), (2739,-0.371645), (2740,-0.422219), (2741,-0.273058), (2742,-0.443468), (2743,-0.480109), (2744,-0.674677), (2745,-0.030361), (2746,-0.199844), (2747,-0.239273), (2748,-0.404579), (2749,-0.409167), (2750,-0.580973), (2751,-0.637584), (2752,-0.805207), (2753,-0.162288), (2754,-0.302510), (2755,-0.337292), (2756,-0.477978), (2757,-0.247064), (2758,-0.391933), (2759,-0.424392), (2760,-0.589228), (2761,0.096420), (2762,-0.088855), (2763,-0.142679), (2764,-0.279645), (2765,-0.302348), (2766,-0.468581), (2767,-0.494540), (2768,-0.683528), (2769,-0.032714), (2770,-0.159930), (2771,-0.201682), (2772,-0.333538), (2773,-0.112850), (2774,-0.281400), (2775,-0.303177), (2776,-0.716520), (2777,-0.044804), (2778,-0.227293), (2779,-0.272757), (2780,-0.427844), (2781,-0.446365), (2782,-0.587514), (2783,-0.644124), (2784,-0.828472), (2785,-0.132605), (2786,-0.313697), (2787,-0.371703), (2788,-0.522144), (2789,-0.278689), (2790,-0.448178), (2791,-0.493636), (2792,-0.546070), (2793,-0.321199), (2794,-0.043373), (2795,-0.203101), (2796,-0.268076), (2797,-0.429200), (2798,-0.422636), (2799,-0.593979), (2800,-0.627834), (2801,-0.388561), (2802,-0.099590), (2803,-0.275572), (2804,-0.321037), (2805,-0.371147), (2806,-0.214554), (2807,-0.374287), (2808,-0.585573), (2809,0.150244), (2810,0.006772), (2811,-0.050771), (2812,-0.236973), (2813,-0.245744), (2814,-0.394789), (2815,-0.450009), (2816,-0.658508), (2817,0.000666), (2818,-0.133984), (2819,-0.207776), (2820,-0.368899), (2821,-0.125450), (2822,-0.262416), (2823,-0.327392), (2824,-0.523349), (2825,-0.280827), (2826,-0.037841), (2827,-0.209647), (2828,-0.264867), (2829,-0.455715), (2830,-0.437542), (2831,-0.589373), (2832,-0.603254), (2833,-0.363055), (2834,-0.088478), (2835,-0.244493), (2836,-0.315968), (2837,-0.418564), (2838,-0.228063), (2839,-0.410088), (2840,-0.187077), (2841,-0.359347), (2842,0.015090), (2843,-0.119089), (2844,-0.128787), (2845,-0.298270), (2846,-0.359526), (2847,-0.493243), (2848,-0.227496), (2849,-0.393266), (2850,-0.070850), (2851,-0.184592), (2852,-0.007567), (2853,-0.175653), (2854,-0.136115), (2855,-0.307921), (2856,-0.638586), (2857,0.030344), (2858,-0.107092), (2859,-0.201792), (2860,-0.374988), (2861,-0.360998), (2862,-0.540237), (2863,-0.589414), (2864,-0.740782), (2865,-0.060243), (2866,-0.213008), (2867,-0.248253), (2868,-0.425632), (2869,-0.178000), (2870,-0.308930), (2871,-0.386441), (2872,-0.316710), (2873,-0.063041), (2874,-0.126621), (2875,-0.313755), (2876,-0.302552), (2877,-0.459956), (2878,-0.517499), (2879,-0.682336), (2880,-0.382212), (2881,-0.109966), (2882,-0.198629), (2883,-0.351851), (2884,-0.193867), (2885,-0.249087), (2886,-0.314520), (2887,-0.477503), (2888,-0.626548), (2889,0.056777), (2890,-0.079726), (2891,-0.172566), (2892,-0.325793), (2893,-0.335491), (2894,-0.462708), (2895,-0.533720), (2896,-0.685088), (2897,-0.005476), (2898,-0.149411), (2899,-0.189302), (2900,-0.362035), (2901,-0.123226), (2902,-0.295502), (2903,-0.349789), (2904,-0.136990), (2905,-0.276749), (2906,0.073537), (2907,-0.056930), (2908,-0.046189), (2909,-0.167364), (2910,-0.248131), (2911,-0.420401), (2912,-0.132819), (2913,-0.315778), (2914,0.001991), (2915,-0.131725), (2916,0.034161), (2917,-0.129286), (2918,-0.099504), (2919,-0.267127), (2920,-0.288903), (2921,-0.007828), (2922,-0.158269), (2923,-0.182362), (2924,-0.407123), (2925,-0.388024), (2926,-0.566329), (2927,-0.646634), (2928,-0.377167), (2929,-0.067757), (2930,-0.227485), (2931,-0.272486), (2932,-0.342101), (2933,-0.214311), (2934,-0.389831), (2935,-0.388846), (2936,-0.587596), (2937,0.092949), (2938,-0.065388), (2939,-0.091804), (2940,-0.275689), (2941,-0.288173), (2942,-0.468808), (2943,-0.514273), (2944,-0.774331), (2945,-0.490932), (2946,-0.248410), (2947,-0.312452), (2948,-0.505160), (2949,-0.331384), (2950,-0.421901), (2951,-0.466902), (2952,-0.820792), (2953,-0.112376), (2954,-0.281395), (2955,-0.357517), (2956,-0.506098), (2957,-0.483286), (2958,-0.650446), (2959,-0.694050), (2960,-0.867716), (2961,-0.195536), (2962,-0.378952), (2963,-0.427202), (2964,-0.592039), (2965,-0.358346), (2966,-0.491135), (2967,-0.548209), (2968,-0.575558), (2969,-0.727389), (2970,-0.059856), (2971,-0.233515), (2972,-0.252505), (2973,-0.432671), (2974,-0.423327), (2975,-0.579341), (2976,-0.648957), (2977,-0.776637), (2978,-0.094238), (2979,-0.272080), (2980,-0.307789), (2981,-0.440579), (2982,-0.222207), (2983,-0.372185), (2984,-0.666620), (2985,-0.469614), (2986,-0.202007), (2987,-0.338979), (2988,-0.360756), (2989,-0.548354), (2990,-0.547369), (2991,-0.702450), (2992,-0.751628), (2993,-0.507715), (2994,-0.215487), (2995,-0.374758), (2996,-0.407210), (2997,-0.533037), (2998,-0.358792), (2999,-0.527348), (3000,-0.605323), (3001,-0.761801), (3002,-0.107272), (3003,-0.257250), (3004,-0.288776), (3005,-0.458723), (3006,-0.448915), (3007,-0.609106), (3008,-0.691733), (3009,-0.841705), (3010,-0.157916), (3011,-0.320430), (3012,-0.348243), (3013,-0.498214), (3014,-0.279849), (3015,-0.402883), (3016,-0.641577), (3017,-0.407413), (3018,-0.124015), (3019,-0.308826), (3020,-0.355217), (3021,-0.529347), (3022,-0.495851), (3023,-0.667657), (3024,-0.733553), (3025,-0.506823), (3026,-0.217851), (3027,-0.389194), (3028,-0.430012), (3029,-0.509847), (3030,-0.347687), (3031,-0.518560), (3032,-0.592358), (3033,-0.724221), (3034,-0.070620), (3035,-0.224774), (3036,-0.287427), (3037,-0.407668), (3038,-0.403434), (3039,-0.552479), (3040,-0.628137), (3041,-0.772999), (3042,-0.096173), (3043,-0.267979), (3044,-0.297188), (3045,-0.400717), (3046,-0.176773), (3047,-0.327208), (3048,-0.370349), (3049,-0.576532), (3050,0.099367), (3051,-0.032026), (3052,-0.093752), (3053,-0.264625), (3054,-0.309163), (3055,-0.442416), (3056,-0.486484), (3057,-0.626706), (3058,0.034791), (3059,-0.104967), (3060,-0.218709), (3061,-0.382619), (3062,-0.113153), (3063,-0.253838), (3064,-0.350861), (3065,-0.520344), (3066,0.125824), (3067,0.016259), (3068,-0.051503), (3069,-0.209370), (3070,-0.234397), (3071,-0.385765), (3072,-0.440521), (3073,-0.625333), (3074,0.066821), (3075,-0.069681), (3076,-0.141626), (3077,-0.279056), (3078,-0.054185), (3079,-0.211126), (3080,-0.429381), (3081,-0.594224), (3082,0.098863), (3083,-0.031140), (3084,-0.097969), (3085,-0.261879), (3086,-0.282259), (3087,-0.419232), (3088,-0.478165), (3089,-0.617924), (3090,0.082126), (3091,-0.104075), (3092,-0.180660), (3093,-0.350143), (3094,-0.118773), (3095,-0.264561), (3096,-0.679302), (3097,-0.395440), (3098,-0.154307), (3099,-0.179797), (3100,-0.315373), (3101,-0.338546), (3102,-0.492231), (3103,-0.547451), (3104,-0.689996), (3105,-0.400091), (3106,-0.165934), (3107,-0.232764), (3108,-0.386918), (3109,-0.255872), (3110,-0.321775), (3111,-0.372812), (3112,-0.562733), (3113,-0.279798), (3114,-0.007551), (3115,-0.078093), (3116,-0.217389), (3117,-0.210361), (3118,-0.387740), (3119,-0.427169), (3120,-0.569714), (3121,-0.294675), (3122,-0.056798), (3123,-0.096683), (3124,-0.291251), (3125,-0.142559), (3126,-0.229827), (3127,-0.288760), (3128,-0.576225), (3129,-0.317911), (3130,-0.054950), (3131,-0.094372), (3132,-0.242027), (3133,-0.223391), (3134,-0.422598), (3135,-0.463416), (3136,-0.636155), (3137,-0.364365), (3138,-0.071681), (3139,-0.111572), (3140,-0.273159), (3141,-0.127248), (3142,-0.187578), (3143,-0.259980), (3144,-0.473589), (3145,-0.213414), (3146,0.038394), (3147,0.021264), (3148,-0.155652), (3149,-0.132369), (3150,-0.339942), (3151,-0.389583), (3152,-0.555353), (3153,-0.266381), (3154,-0.014566), (3155,-0.076286), (3156,-0.235087), (3157,-0.093828), (3158,-0.184808), (3159,-0.250711), (3160,-0.614356), (3161,-0.367650), (3162,-0.120018), (3163,-0.176165), (3164,-0.329393), (3165,-0.293105), (3166,-0.483489), (3167,-0.520594), (3168,-0.677999), (3169,-0.399246), (3170,-0.144645), (3171,-0.207761), (3172,-0.364702), (3173,-0.204858), (3174,-0.280053), (3175,-0.346882), (3176,-0.732355), (3177,-0.043914), (3178,-0.195752), (3179,-0.248649), (3180,-0.393048), (3181,-0.407855), (3182,-0.545291), (3183,-0.617693), (3184,-0.756982), (3185,-0.064364), (3186,-0.218518), (3187,-0.271879), (3188,-0.437649), (3189,-0.197913), (3190,-0.322343), (3191,-0.397995), (3192,-0.589312), (3193,-0.328205), (3194,-0.094048), (3195,-0.162737), (3196,-0.335470), (3197,-0.322870), (3198,-0.442654), (3199,-0.511343), (3200,-0.839221), (3201,-0.593912), (3202,-0.364395), (3203,-0.422859), (3204,-0.559368), (3205,-0.442724), (3206,-0.514199), (3207,-0.518787), (3208,-0.858738), (3209,-0.222788), (3210,-0.367657), (3211,-0.436339), (3212,-0.603969), (3213,-0.603911), (3214,-0.739024), (3215,-0.803066), (3216,-0.949325), (3217,-0.279468), (3218,-0.434549), (3219,-0.511598), (3220,-0.648570), (3221,-0.431132), (3222,-0.580640), (3223,-0.613562), (3224,-0.636266), (3225,-0.773232), (3226,-0.098266), (3227,-0.244524), (3228,-0.348053), (3229,-0.505457), (3230,-0.498899), (3231,-0.667919), (3232,-0.744504), (3233,-0.889836), (3234,-0.247380), (3235,-0.357409), (3236,-0.452109), (3237,-0.601617), (3238,-0.361881), (3239,-0.490957), (3240,-0.813256), (3241,-0.560515), (3242,-0.306383), (3243,-0.445672), (3244,-0.492997), (3245,-0.678735), (3246,-0.672177), (3247,-0.837014), (3248,-0.885265), (3249,-0.621841), (3250,-0.317077), (3251,-0.448934), (3252,-0.549670), (3253,-0.598854), (3254,-0.467345), (3255,-0.653546), (3256,-0.711089), (3257,-0.861531), (3258,-0.169840), (3259,-0.368590), (3260,-0.385250), (3261,-0.538015), (3262,-0.577437), (3263,-0.759462), (3264,-0.794244), (3265,-0.954904), (3266,-0.278078), (3267,-0.414118), (3268,-0.459582), (3269,-0.603981), (3270,-0.394438), (3271,-0.504004), (3272,-0.727368), (3273,-0.505747), (3274,-0.231641), (3275,-0.373253), (3276,-0.437759), (3277,-0.603066), (3278,-0.609044), (3279,-0.783637), (3280,-0.838393), (3281,-0.580079), (3282,-0.292497), (3283,-0.457797), (3284,-0.511158), (3285,-0.548726), (3286,-0.435802), (3287,-0.618290), (3288,-0.681400), (3289,-0.835561), (3290,-0.150369), (3291,-0.282695), (3292,-0.330946), (3293,-0.499039), (3294,-0.514773), (3295,-0.679610), (3296,-0.758518), (3297,-0.920568), (3298,-0.234920), (3299,-0.399756), (3300,-0.451263), (3301,-0.624923), (3302,-0.432569), (3303,-0.555140), (3304,-0.580629), (3305,-0.739430), (3306,-0.103943), (3307,-0.260884), (3308,-0.320281), (3309,-0.427523), (3310,-0.442330), (3311,-0.576046), (3312,-0.622907), (3313,-0.773349), (3314,-0.107668), (3315,-0.253464), (3316,-0.297068), (3317,-0.459119), (3318,-0.218456), (3319,-0.369824), (3320,-0.523978), (3321,-0.692998), (3322,-0.008276), (3323,-0.163827), (3324,-0.254807), (3325,-0.410822), (3326,-0.411697), (3327,-0.589076), (3328,-0.689348), (3329,-0.777549), (3330,-0.091430), (3331,-0.247445), (3332,-0.324029), (3333,-0.468428), (3334,-0.252386), (3335,-0.380993), (3336,-0.607144), (3337,-0.758976), (3338,-0.080296), (3339,-0.249316), (3340,-0.307316), (3341,-0.470300), (3342,-0.489753), (3343,-0.624396), (3344,-0.692622), (3345,-0.851886), (3346,-0.182492), (3347,-0.337110), (3348,-0.377002), (3349,-0.492603), (3350,-0.283061), (3351,-0.454867), (3352,-0.727467), (3353,-0.451501), (3354,-0.223844), (3355,-0.250730), (3356,-0.423926), (3357,-0.400180), (3358,-0.576169), (3359,-0.618847), (3360,-0.816664), (3361,-0.548594), (3362,-0.290273), (3363,-0.323665), (3364,-0.495001), (3365,-0.344450), (3366,-0.425681), (3367,-0.509699), (3368,-0.683365), (3369,-0.409252), (3370,-0.133749), (3371,-0.184786), (3372,-0.347770), (3373,-0.352358), (3374,-0.545066), (3375,-0.610968), (3376,-0.734002), (3377,-0.450603), (3378,-0.180210), (3379,-0.250295), (3380,-0.422565), (3381,-0.286873), (3382,-0.339770), (3383,-0.415428), (3384,-0.793932), (3385,-0.531898), (3386,-0.314923), (3387,-0.348308), (3388,-0.477848), (3389,-0.457815), (3390,-0.619409), (3391,-0.688091), (3392,-0.858044), (3393,-0.565816), (3394,-0.322831), (3395,-0.336711), (3396,-0.496438), (3397,-0.342631), (3398,-0.441514), (3399,-0.485119), (3400,-0.741927), (3401,-0.436700), (3402,-0.209969), (3403,-0.273549), (3404,-0.443495), (3405,-0.393738), (3406,-0.583659), (3407,-0.652812), (3408,-0.768413), (3409,-0.485014), (3410,-0.242961), (3411,-0.255446), (3412,-0.448616), (3413,-0.298992), (3414,-0.397875), (3415,-0.474923), (3416,-0.738701), (3417,-0.446936), (3418,-0.207670), (3419,-0.250341), (3420,-0.397070), (3421,-0.428132), (3422,-0.597615), (3423,-0.636110), (3424,-0.775406), (3425,-0.494794), (3426,-0.223004), (3427,-0.267542), (3428,-0.425409), (3429,-0.285077), (3430,-0.372808), (3431,-0.406200), (3432,-0.791203), (3433,-0.146894), (3434,-0.293616), (3435,-0.342337), (3436,-0.504850), (3437,-0.519194), (3438,-0.642691), (3439,-0.728099), (3440,-0.905015), (3441,-0.237018), (3442,-0.395355), (3443,-0.431064), (3444,-0.569426), (3445,-0.339909), (3446,-0.526580), (3447,-0.585514), (3448,-0.748027), (3449,-0.493896), (3450,-0.234648), (3451,-0.269894), (3452,-0.456565), (3453,-0.413771), (3454,-0.605552), (3455,-0.643584), (3456,-1.011405), (3457,-0.717787), (3458,-0.457150), (3459,-0.524449), (3460,-0.671171), (3461,-0.532229), (3462,-0.571657), (3463,-0.598536), (3464,-0.759660), (3465,-0.463719), (3466,-0.231416), (3467,-0.263411), (3468,-0.415706), (3469,-0.408685), (3470,-0.606502), (3471,-0.687263), (3472,-0.825163), (3473,-0.563135), (3474,-0.318290), (3475,-0.347492), (3476,-0.523018), (3477,-0.387789), (3478,-0.506183), (3479,-0.553038), (3480,-0.840503), (3481,-0.967256), (3482,-0.287174), (3483,-0.447371), (3484,-0.522097), (3485,-0.645594), (3486,-0.666907), (3487,-0.794124), (3488,-0.886031), (3489,-1.040655), (3490,-0.368475), (3491,-0.490113), (3492,-0.530004), (3493,-0.685085), (3494,-0.467647), (3495,-0.609260), (3496,-0.713252), (3497,-0.882271), (3498,-0.197550), (3499,-0.323833), (3500,-0.366048), (3501,-0.510447), (3502,-0.509462), (3503,-0.688701), (3504,-0.754603), (3505,-0.925476), (3506,-0.232858), (3507,-0.401415), (3508,-0.476140), (3509,-0.631691), (3510,-0.381272), (3511,-0.554938), (3512,-0.867951), (3513,-1.029075), (3514,-0.357822), (3515,-0.491538), (3516,-0.533283), (3517,-0.677225), (3518,-0.695282), (3519,-0.853149), (3520,-0.936240), (3521,-1.068097), (3522,-0.401490), (3523,-0.542645), (3524,-0.574171), (3525,-0.719966), (3526,-0.470474), (3527,-0.645530), (3528,-0.662661), (3529,-0.828894), (3530,-0.156714), (3531,-0.278358), (3532,-0.285733), (3533,-0.445460), (3534,-0.463517), (3535,-0.628354), (3536,-0.664069), (3537,-0.835405), (3538,-0.201315), (3539,-0.358256), (3540,-0.393501), (3541,-0.570880), (3542,-0.321395), (3543,-0.454185), (3544,-0.786240), (3545,-0.898128), (3546,-0.219905), (3547,-0.382419), (3548,-0.462260), (3549,-0.631280), (3550,-0.656769), (3551,-0.790022), (3552,-0.829914), (3553,-1.006360), (3554,-0.336503), (3555,-0.485085), (3556,-0.544481), (3557,-0.658693), (3558,-0.435682), (3559,-0.571721), (3560,-0.602320), (3561,-0.770876), (3562,-0.096374), (3563,-0.257491), (3564,-0.303419), (3565,-0.458043), (3566,-0.457522), (3567,-0.616322), (3568,-0.696620), (3569,-0.852634), (3570,-0.183704), (3571,-0.330426), (3572,-0.381000), (3573,-0.514723), (3574,-0.268944), (3575,-0.465371), (3576,-0.428156), (3577,-0.578591), (3578,-0.286370), (3579,-0.021086), (3580,-0.067014), (3581,-0.213736), (3582,-0.228543), (3583,-0.419397), (3584,-0.515024), (3585,-0.682647), (3586,-0.380670), (3587,-0.138148), (3588,-0.217982), (3589,-0.356345), (3590,-0.189538), (3591,-0.270300), (3592,-0.479269), (3593,-0.654325), (3594,-0.352348), (3595,-0.130727), (3596,-0.152503), (3597,-0.320590), (3598,-0.305210), (3599,-0.506740), (3600,-0.562887), (3601,-0.704499), (3602,-0.394626), (3603,-0.153963), (3604,-0.244017), (3605,-0.396311), (3606,-0.233218), (3607,-0.287512), (3608,-0.544783), (3609,-0.288792), (3610,-0.447593), (3611,-0.136786), (3612,-0.286758), (3613,-0.271841), (3614,-0.450617), (3615,-0.513726), (3616,-0.650235), (3617,-0.365440), (3618,-0.534460), (3619,-0.173492), (3620,-0.309068), (3621,-0.169199), (3622,-0.340542), (3623,-0.326545), (3624,-0.748718), (3625,-0.441162), (3626,-0.228370), (3627,-0.281730), (3628,-0.428452), (3629,-0.424681), (3630,-0.558397), (3631,-0.614544), (3632,-0.788210), (3633,-0.521993), (3634,-0.270185), (3635,-0.309606), (3636,-0.471663), (3637,-0.332258), (3638,-0.411159), (3639,-0.453837), (3640,-0.582444), (3641,-0.287900), (3642,-0.441591), (3643,-0.125212), (3644,-0.304451), (3645,-0.319721), (3646,-0.463193), (3647,-0.532352), (3648,-0.711584), (3649,-0.492756), (3650,-0.632508), (3651,-0.272467), (3652,-0.414085), (3653,-0.256095), (3654,-0.372166), (3655,-0.356780), (3656,-0.624734), (3657,-0.342732), (3658,-0.473662), (3659,-0.124772), (3660,-0.284036), (3661,-0.281655), (3662,-0.416768), (3663,-0.460372), (3664,-0.629855), (3665,-0.338097), (3666,-0.510367), (3667,-0.156831), (3668,-0.274755), (3669,-0.147429), (3670,-0.315052), (3671,-0.262972), (3672,-0.523030), (3673,-0.277721), (3674,-0.422126), (3675,-0.089956), (3676,-0.224599), (3677,-0.218504), (3678,-0.384274), (3679,-0.446457), (3680,-0.616873), (3681,-0.333475), (3682,-0.496915), (3683,-0.163817), (3684,-0.304966), (3685,-0.164634), (3686,-0.332721), (3687,-0.298756), (3688,-0.684699), (3689,-0.423128), (3690,-0.211726), (3691,-0.249758), (3692,-0.409955), (3693,-0.407574), (3694,-0.583093), (3695,-0.649929), (3696,-0.795254), (3697,-0.493277), (3698,-0.227993), (3699,-0.282287), (3700,-0.481031), (3701,-0.300286), (3702,-0.363402), (3703,-0.404683), (3704,-0.793406), (3705,-0.503045), (3706,-0.307435), (3707,-0.340820), (3708,-0.493585), (3709,-0.488417), (3710,-0.644431), (3711,-0.695932), (3712,-0.760901), (3713,-0.923421), (3714,-0.234517), (3715,-0.410506), (3716,-0.449464), (3717,-0.618484), (3718,-0.356456), (3719,-0.505038), (3720,-0.828733), (3721,-0.590850), (3722,-0.274478), (3723,-0.426309), (3724,-0.505217), (3725,-0.657975), (3726,-0.667210), (3727,-0.813468), (3728,-0.836171), (3729,-0.608514), (3730,-0.324189), (3731,-0.480196), (3732,-0.543312), (3733,-0.605502), (3734,-0.499070), (3735,-0.625360), (3736,-0.646204), (3737,-0.740904), (3738,-0.489559), (3739,-0.212196), (3740,-0.358455), (3741,-0.437362), (3742,-0.583621), (3743,-0.585886), (3744,-0.731681), (3745,-0.810126), (3746,-0.556451), (3747,-0.278632), (3748,-0.438822), (3749,-0.502865), (3750,-0.567377), (3751,-0.405211), (3752,-0.816695), (3753,-0.477092), (3754,-0.651684), (3755,-0.358530), (3756,-0.524763), (3757,-0.595312), (3758,-0.729491), (3759,-0.685771), (3760,-0.841785), (3761,-0.486389), (3762,-0.634508), (3763,-0.399418), (3764,-0.552646), (3765,-0.539119), (3766,-0.694663), (3767,-0.508345), (3768,-0.681548), (3769,-0.765565), (3770,-0.552767), (3771,-0.240108), (3772,-0.400768), (3773,-0.405819), (3774,-0.606886), (3775,-0.610548), (3776,-0.751697), (3777,-0.793905), (3778,-0.550919), (3779,-0.289355), (3780,-0.455118), (3781,-0.495473), (3782,-0.542334), (3783,-0.395496), (3784,-0.760068), (3785,-0.420464), (3786,-0.582978), (3787,-0.318627), (3788,-0.469532), (3789,-0.569341), (3790,-0.701661), (3791,-0.696500), (3792,-0.837186), (3793,-0.499905), (3794,-0.669852), (3795,-0.385990), (3796,-0.522029), (3797,-0.519648), (3798,-0.681698), (3799,-0.520002), (3800,-0.667650), (3801,-0.710791), (3802,-0.453404), (3803,-0.163505), (3804,-0.320910), (3805,-0.385885), (3806,-0.560941), (3807,-0.562280), (3808,-0.707142), (3809,-0.788836), (3810,-0.540741), (3811,-0.277317), (3812,-0.423112), (3813,-0.478332), (3814,-0.551197), (3815,-0.400646), (3816,-0.561300), (3817,-0.577967), (3818,-0.335908), (3819,-0.090136), (3820,-0.247077), (3821,-0.313906), (3822,-0.463884), (3823,-0.452680), (3824,-0.614731), (3825,-0.678773), (3826,-0.447866), (3827,-0.163534), (3828,-0.345096), (3829,-0.386378), (3830,-0.423483), (3831,-0.295223), (3832,-0.575256), (3833,-0.618867), (3834,-0.370765), (3835,-0.129639), (3836,-0.287043), (3837,-0.311143), (3838,-0.455542), (3839,-0.455953), (3840,-0.631936), (3841,-0.686693), (3842,-0.464139), (3843,-0.197002), (3844,-0.346510), (3845,-0.406376), (3846,-0.429079), (3847,-0.287351), (3848,-0.657032), (3849,-0.717825), (3850,-0.437213), (3851,-0.149168), (3852,-0.313078), (3853,-0.349713), (3854,-0.542421), (3855,-0.527041), (3856,-0.719285), (3857,-0.734092), (3858,-0.515257), (3859,-0.219317), (3860,-0.333991), (3861,-0.414289), (3862,-0.492734), (3863,-0.302697), (3864,-0.616173), (3865,-0.769864), (3866,-0.096758), (3867,-0.215146), (3868,-0.268043), (3869,-0.429166), (3870,-0.443973), (3871,-0.601841), (3872,-0.682609), (3873,-0.854878), (3874,-0.188735), (3875,-0.321988), (3876,-0.405078), (3877,-0.529039), (3878,-0.275834), (3879,-0.421629), (3880,-0.537694), (3881,-0.694172), (3882,-0.002487), (3883,-0.156178), (3884,-0.229970), (3885,-0.408745), (3886,-0.433772), (3887,-0.595822), (3888,-0.618995), (3889,-0.752711), (3890,-0.116298), (3891,-0.281135), (3892,-0.335422), (3893,-0.474718), (3894,-0.231262), (3895,-0.411897), (3896,-0.661273), (3897,-0.790806), (3898,-0.111194), (3899,-0.261172), (3900,-0.327075), (3901,-0.479369), (3902,-0.475598), (3903,-0.640435), (3904,-0.683576), (3905,-0.845163), (3906,-0.179489), (3907,-0.364301), (3908,-0.421375), (3909,-0.585748), (3910,-0.306069), (3911,-0.462083), (3912,-0.633889), (3913,-0.799653), (3914,-0.124687), (3915,-0.301602), (3916,-0.371681), (3917,-0.534201), (3918,-0.555978), (3919,-0.701766), (3920,-0.763492), (3921,-0.914860), (3922,-0.225492), (3923,-0.353173), (3924,-0.420928), (3925,-0.557901), (3926,-0.333957), (3927,-0.475569), (3928,-0.627870), (3929,-0.821041), (3930,-0.128887), (3931,-0.254244), (3932,-0.298781), (3933,-0.446430), (3934,-0.468670), (3935,-0.640476), (3936,-0.707305), (3937,-0.836381), (3938,-0.142367), (3939,-0.308600), (3940,-0.348492), (3941,-0.504969), (3942,-0.289848), (3943,-0.437966), (3944,-0.728218), (3945,-0.516816), (3946,-0.265934), (3947,-0.423802), (3948,-0.418641), (3949,-0.619708), (3950,-0.653093), (3951,-0.814217), (3952,-0.846676), (3953,-0.616695), (3954,-0.330974), (3955,-0.441929), (3956,-0.472528), (3957,-0.544936), (3958,-0.395775), (3959,-0.535997), (3960,-0.584712), (3961,-0.760231), (3962,-0.061113), (3963,-0.222701), (3964,-0.287670), (3965,-0.432538), (3966,-0.470570), (3967,-0.642376), (3968,-0.522013), (3969,-0.267881), (3970,0.027596), (3971,-0.152106), (3972,-0.224977), (3973,-0.273228), (3974,-0.142182), (3975,-0.307952), (3976,-0.407761), (3977,-0.197750), (3978,0.088899), (3979,-0.062006), (3980,-0.092605), (3981,-0.285312), (3982,-0.294547), (3983,-0.468676), (3984,-0.502525), (3985,-0.251180), (3986,0.035006), (3987,-0.141910), (3988,-0.179472), (3989,-0.250948), (3990,-0.096214), (3991,-0.278709), (3992,-0.440759), (3993,-0.113234), (3994,-0.237195), (3995,-0.008605), (3996,-0.175771), (3997,-0.268611), (3998,-0.407437), (3999,-0.391587), (4000,-0.518804), (4001,-0.196852), (4002,-0.303630), (4003,-0.029518), (4004,-0.190641), (4005,-0.184084), (4006,-0.317337), (4007,-0.177005), (4008,-0.221536), (4009,-0.269324), (4010,-0.391431), (4011,-0.092704), (4012,-0.288198), (4013,-0.345271), (4014,-0.536589), (4015,-0.541177), (4016,-0.274966), (4017,-0.339472), (4018,-0.470402), (4019,-0.173998), (4020,-0.231541), (4021,-0.303943), (4022,-0.458561), (4023,-0.317302), (4024,-0.523015), (4025,-0.168083), (4026,-0.304586), (4027,-0.031406), (4028,-0.163733), (4029,-0.239854), (4030,-0.390759), (4031,-0.366080), (4032,-0.529990), (4033,-0.232196), (4034,-0.402606), (4035,-0.113634), (4036,-0.254783), (4037,-0.219428), (4038,-0.356857), (4039,-0.236964), (4040,-0.439427), (4041,-0.073812), (4042,-0.237723), (4043,0.042426), (4044,-0.080144), (4045,-0.179027), (4046,-0.324822), (4047,-0.347055), (4048,-0.483095), (4049,-0.164863), (4050,-0.331096), (4051,-0.031905), (4052,-0.194419), (4053,-0.174392), (4054,-0.319718), (4055,-0.166844), (4056,-0.439444), (4057,-0.106346), (4058,-0.246105), (4059,0.027544), (4060,-0.115928), (4061,-0.145601), (4062,-0.336455), (4063,-0.346616), (4064,-0.495661), (4065,-0.152807), (4066,-0.296743), (4067,-0.044001), (4068,-0.204192), (4069,-0.202280), (4070,-0.341570), (4071,-0.159435), (4072,-0.327058), (4073,0.040416), (4074,-0.160194), (4075,0.133894), (4076,-0.026303), (4077,-0.116357), (4078,-0.229635), (4079,-0.215182), (4080,-0.423218), (4081,-0.060390), (4082,-0.215014), (4083,0.062349), (4084,-0.109921), (4085,-0.073633), (4086,-0.225470), (4087,-0.062371), (4088,-0.371208), (4089,-0.026031), (4090,-0.172290), (4091,0.108323), (4092,-0.034223), (4093,-0.127526), (4094,-0.270535), (4095,-0.288129), (4096,-0.469227), (4097,-0.144482), (4098,-0.273559), (4099,-0.009672), (4100,-0.145711), (4101,-0.125678), (4102,-0.272400), (4103,-0.113490), (4104,-0.414424), (4105,-0.051596), (4106,-0.215043), (4107,0.052101), (4108,-0.117382), (4109,-0.183285), (4110,-0.328617), (4111,-0.293255), (4112,-0.464598), (4113,-0.146829), (4114,-0.265680), (4115,0.001927), (4116,-0.159667), (4117,-0.157286), (4118,-0.284966), (4119,-0.147884), (4120,-0.249546), (4121,-0.398128), (4122,0.243395), (4123,0.072052), (4124,0.003363), (4125,-0.132213), (4126,-0.135405), (4127,-0.301638), (4128,-0.351749), (4129,-0.503580), (4130,0.167673), (4131,0.000043), (4132,-0.062603), (4133,-0.254384), (4134,0.043417), (4135,-0.084733), (4136,-0.295092), (4137,-0.062783), (4138,0.202964), (4139,0.069711), (4140,0.004272), (4141,-0.166137), (4142,-0.168872), (4143,-0.358330), (4144,-0.374990), (4145,-0.143620), (4146,0.139315), (4147,-0.027845), (4148,-0.061230), (4149,-0.102981), (4150,0.054539), (4151,-0.120517), (4152,-0.382435), (4153,-0.130620), (4154,0.149523), (4155,-0.006955), (4156,-0.057059), (4157,-0.195422), (4158,-0.192114), (4159,-0.355561), (4160,-0.421463), (4161,-0.180331), (4162,0.120250), (4163,-0.077567), (4164,-0.090051), (4165,-0.178715), (4166,-0.027694), (4167,-0.189281), (4168,-0.333680), (4169,-0.059574), (4170,0.199668), (4171,0.028794), (4172,-0.013420), (4173,-0.184763), (4174,-0.176809), (4175,-0.367657), (4176,-0.402439), (4177,-0.164562), (4178,0.117446), (4179,-0.032068), (4180,-0.082636), (4181,-0.164330), (4182,-0.010993), (4183,-0.179549), (4184,-0.238946), (4185,-0.387527), (4186,0.271184), (4187,0.096591), (4188,0.053913), (4189,-0.087236), (4190,-0.102976), (4191,-0.236229), (4192,-0.297485), (4193,-0.421909), (4194,0.245624), (4195,0.106335), (4196,0.015812), (4197,-0.130910), (4198,0.094424), (4199,-0.070413), (4200,-0.050380), (4201,-0.198962), (4202,0.074218), (4203,-0.070187), (4204,-0.132370), (4205,-0.306036), (4206,-0.279034), (4207,-0.444340), (4208,-0.088482), (4209,-0.238923), (4210,0.022648), (4211,-0.136153), (4212,-0.069671), (4213,-0.238691), (4214,-0.114614), (4215,-0.237648), (4216,-0.358359), (4217,-0.126988), (4218,0.131326), (4219,-0.000067), (4220,-0.045068), (4221,-0.230343), (4222,-0.195445), (4223,-0.373757), (4224,-0.430367), (4225,-0.176699), (4226,-0.086066), (4227,-0.233715), (4228,-0.281965), (4229,-0.373415), (4230,-0.090017), (4231,-0.227452), (4232,-0.383467), (4233,-0.152553), (4234,-0.129740), (4235,-0.290394), (4236,-0.314494), (4237,-0.484440), (4238,-0.197792), (4239,-0.380280), (4240,-0.402520), (4241,-0.160461), (4242,-0.029878), (4243,-0.181716), (4244,-0.221601), (4245,-0.262889), (4246,-0.008288), (4247,-0.178698), (4248,-0.468486), (4249,-0.224574), (4250,-0.231015), (4251,-0.355909), (4252,-0.406946), (4253,-0.604763), (4254,-0.303249), (4255,-0.461587), (4256,-0.526562), (4257,-0.270101), (4258,-0.123263), (4259,-0.286710), (4260,-0.338211), (4261,-0.399467), (4262,-0.105386), (4263,-0.269296), (4264,-0.323583), (4265,0.019733), (4266,-0.147896), (4267,-0.152484), (4268,-0.318711), (4269,-0.384150), (4270,-0.535982), (4271,-0.292069), (4272,-0.445760), (4273,-0.122875), (4274,-0.265884), (4275,-0.110687), (4276,-0.257872), (4277,-0.222054), (4278,-0.425444), (4279,-0.132289), (4280,-0.433693), (4281,-0.219505), (4282,-0.206441), (4283,-0.308110), (4284,-0.378189), (4285,-0.560215), (4286,-0.248945), (4287,-0.416105), (4288,-0.477361), (4289,-0.265959), (4290,-0.086611), (4291,-0.254234), (4292,-0.271364), (4293,-0.358168), (4294,-0.080812), (4295,-0.239606), (4296,-0.350105), (4297,0.002041), (4298,-0.131675), (4299,-0.117685), (4300,-0.273699), (4301,-0.348888), (4302,-0.501652), (4303,-0.225223), (4304,-0.373335), (4305,-0.028158), (4306,-0.170704), (4307,-0.039194), (4308,-0.182666), (4309,-0.125013), (4310,-0.287064), (4311,-0.042218), (4312,-0.402144), (4313,-0.155908), (4314,-0.190220), (4315,-0.371782), (4316,-0.401918), (4317,-0.593699), (4318,-0.279180), (4319,-0.459808), (4320,-0.519675), (4321,-0.257177), (4322,-0.124741), (4323,-0.265427), (4324,-0.311818), (4325,-0.394439), (4326,-0.128229), (4327,-0.268451), (4328,-0.325524), (4329,0.017792), (4330,-0.140545), (4331,-0.142810), (4332,-0.298824), (4333,-0.367044), (4334,-0.504479), (4335,-0.252201), (4336,-0.387777), (4337,-0.026809), (4338,-0.180500), (4339,-0.041095), (4340,-0.225443), (4341,-0.188228), (4342,-0.351669), (4343,-0.068270), (4344,-0.143001), (4345,-0.294369), (4346,0.120481), (4347,-0.048533), (4348,-0.100040), (4349,-0.215641), (4350,0.023168), (4351,-0.140279), (4352,-0.258666), (4353,-0.397962), (4354,0.180856), (4355,-0.001632), (4356,-0.057779), (4357,-0.195678), (4358,0.166687), (4359,-0.004656), (4360,-0.224771), (4361,-0.283241), (4362,-0.052328), (4363,-0.019759), (4364,-0.218966), (4365,-0.244925), (4366,-0.423694), (4367,-0.132869), (4368,-0.285628), (4369,-0.356176), (4370,-0.135018), (4371,0.047116), (4372,-0.100532), (4373,-0.141350), (4374,-0.254165), (4375,0.068250), (4376,-0.221539), (4377,-0.399381), (4378,0.000141), (4379,-0.134972), (4380,-0.165571), (4381,-0.299288), (4382,-0.057698), (4383,-0.212779), (4384,-0.269389), (4385,-0.419831), (4386,0.140872), (4387,-0.020715), (4388,-0.096373), (4389,-0.241241), (4390,0.112764), (4391,-0.035817), (4392,-0.374378), (4393,-0.123496), (4394,-0.089531), (4395,-0.239503), (4396,-0.291473), (4397,-0.491144), (4398,-0.211465), (4399,-0.360973), (4400,-0.385536), (4401,-0.152769), (4402,-0.013827), (4403,-0.205145), (4404,-0.238067), (4405,-0.317901), (4406,-0.041472), (4407,-0.210022), (4408,-0.237835), (4409,-0.343223), (4410,0.055372), (4411,-0.102033), (4412,-0.179081), (4413,-0.286786), (4414,-0.034045), (4415,-0.193778), (4416,-0.267107), (4417,-0.398507), (4418,0.145941), (4419,-0.037017), (4420,-0.081548), (4421,-0.213875), (4422,0.161032), (4423,-0.008921), (4424,-0.182117), (4425,-0.351136), (4426,0.060927), (4427,-0.131317), (4428,-0.149374), (4429,-0.303998), (4430,-0.063792), (4431,-0.207734), (4432,-0.270380), (4433,-0.412462), (4434,0.143595), (4435,-0.038431), (4436,-0.087145), (4437,-0.255231), (4438,0.119669), (4439,-0.022407), (4440,-0.171452), (4441,-0.333045), (4442,0.062300), (4443,-0.083032), (4444,-0.133606), (4445,-0.289150), (4446,-0.037342), (4447,-0.189173), (4448,-0.262508), (4449,-0.412480), (4450,0.139394), (4451,-0.027765), (4452,-0.056975), (4453,-0.201373), (4454,0.148449), (4455,0.001258), (4456,-0.263447), (4457,-0.026497), (4458,-0.017616), (4459,-0.161552), (4460,-0.215375), (4461,-0.384395), (4462,-0.107966), (4463,-0.221707), (4464,-0.234191), (4465,-0.025576), (4466,0.132408), (4467,-0.035215), (4468,-0.086253), (4469,-0.163770), (4470,0.120561), (4471,-0.034526), (4472,-0.265323), (4473,-0.025124), (4474,-0.024603), (4475,-0.178757), (4476,-0.249769), (4477,-0.394631), (4478,-0.120525), (4479,-0.277466), (4480,-0.520342), (4481,-0.241589), (4482,-0.104037), (4483,-0.283740), (4484,-0.325954), (4485,-0.390930), (4486,-0.099165), (4487,-0.271441), (4488,-0.329441), (4489,-0.009349), (4490,-0.161650), (4491,-0.146264), (4492,-0.308778), (4493,-0.387686), (4494,-0.534877), (4495,-0.244509), (4496,-0.384262), (4497,-0.039555), (4498,-0.183490), (4499,-0.038512), (4500,-0.171295), (4501,-0.160092), (4502,-0.305887), (4503,-0.072657), (4504,-0.432582), (4505,-0.080900), (4506,-0.229482), (4507,-0.234539), (4508,-0.400766), (4509,-0.466669), (4510,-0.602245), (4511,-0.332315), (4512,-0.507841), (4513,-0.156158), (4514,-0.334934), (4515,-0.194138), (4516,-0.363621), (4517,-0.340802), (4518,-0.492633), (4519,-0.204125), (4520,-0.374078), (4521,-0.036798), (4522,-0.173764), (4523,-0.163956), (4524,-0.357127), (4525,-0.412347), (4526,-0.552100), (4527,-0.267774), (4528,-0.434934), (4529,-0.052601), (4530,-0.223474), (4531,-0.080819), (4532,-0.223828), (4533,-0.235849), (4534,-0.376065), (4535,-0.104745), (4536,-0.502297), (4537,-0.136219), (4538,-0.302452), (4539,-0.297748), (4540,-0.458872), (4541,-0.526634), (4542,-0.707263), (4543,-0.430833), (4544,-0.615181), (4545,-0.241671), (4546,-0.375851), (4547,-0.256420), (4548,-0.395709), (4549,-0.364067), (4550,-0.521941), (4551,-0.257121), (4552,-0.372259), (4553,-0.036838), (4554,-0.168232), (4555,-0.143559), (4556,-0.276342), (4557,-0.345964), (4558,-0.495472), (4559,-0.252950), (4560,-0.436835), (4561,-0.139034), (4562,-0.291335), (4563,-0.154253), (4564,-0.299579), (4565,-0.276766), (4566,-0.394690), (4567,-0.099213), (4568,-0.552036), (4569,-0.200360), (4570,-0.340576), (4571,-0.346097), (4572,-0.499325), (4573,-0.575440), (4574,-0.706840), (4575,-0.389065), (4576,-0.552511), (4577,-0.187360), (4578,-0.313650), (4579,-0.212335), (4580,-0.344191), (4581,-0.350176), (4582,-0.475996), (4583,-0.187951), (4584,-0.330960), (4585,0.021649), (4586,-0.150157), (4587,-0.145923), (4588,-0.260591), (4589,-0.354364), (4590,-0.534993), (4591,-0.257637), (4592,-0.418761), (4593,-0.081944), (4594,-0.229129), (4595,-0.073931), (4596,-0.233195), (4597,-0.191804), (4598,-0.348282), (4599,-0.102966), (4600,-0.156796), (4601,-0.237094), (4602,-0.016400), (4603,0.012455), (4604,-0.171893), (4605,-0.183914), (4606,-0.344111), (4607,-0.093223), (4608,-0.222762), (4609,-0.294701), (4610,-0.016875), (4611,0.103945), (4612,-0.063678), (4613,-0.099387), (4614,-0.159716), (4615,0.085129), (4616,-0.204659), (4617,-0.269629), (4618,-0.030356), (4619,-0.026121), (4620,-0.183526), (4621,-0.239672), (4622,-0.443069), (4623,-0.143878), (4624,-0.307318), (4625,-0.327235), (4626,-0.084249), (4627,0.082094), (4628,-0.072524), (4629,-0.141676), (4630,-0.192250), (4631,0.117159), (4632,-0.233010), (4633,-0.390884), (4634,0.022576), (4635,-0.125079), (4636,-0.195158), (4637,-0.354892), (4638,-0.091931), (4639,-0.244689), (4640,-0.310592), (4641,-0.452667), (4642,0.083878), (4643,-0.081428), (4644,-0.137105), (4645,-0.295443), (4646,0.119871), (4647,-0.047289), (4648,-0.351943), (4649,-0.090373), (4650,-0.044335), (4651,-0.249122), (4652,-0.285757), (4653,-0.495653), (4654,-0.172305), (4655,-0.354330), (4656,-0.398404), (4657,-0.168417), (4658,-0.036445), (4659,-0.206861), (4660,-0.254178), (4661,-0.342379), (4662,-0.072912), (4663,-0.226140), (4664,-0.283683), (4665,-0.426692), (4666,-0.025774), (4667,-0.132553), (4668,-0.197985), (4669,-0.323806), (4670,-0.071064), (4671,-0.236834), (4672,-0.306450), (4673,-0.426234), (4674,0.124714), (4675,-0.037807), (4676,-0.058650), (4677,-0.211878), (4678,0.140268), (4679,-0.018069), (4680,-0.181046), (4681,-0.307337), (4682,0.075930), (4683,-0.047104), (4684,-0.105111), (4685,-0.269948), (4686,-0.018603), (4687,-0.187153), (4688,-0.252128), (4689,-0.383985), (4690,0.166030), (4691,-0.008563), (4692,-0.076319), (4693,-0.220254), (4694,0.153720), (4695,0.013034), (4696,-0.155059), (4697,-0.332438), (4698,0.074516), (4699,-0.078712), (4700,-0.123243), (4701,-0.316420), (4702,-0.085044), (4703,-0.219687), (4704,-0.234030), (4705,-0.388185), (4706,0.136752), (4707,-0.036451), (4708,-0.090738), (4709,-0.228174), (4710,0.119789), (4711,-0.048298), (4712,-0.285138), (4713,0.073044), (4714,-0.101548), (4715,-0.107996), (4716,-0.252858), (4717,-0.327120), (4718,-0.419497), (4719,-0.138884), (4720,-0.309764), (4721,0.040059), (4722,-0.121065), (4723,0.026700), (4724,-0.081006), (4725,-0.051687), (4726,-0.216524), (4727,0.056656), (4728,-0.349255), (4729,-0.121598), (4730,-0.117827), (4731,-0.278951), (4732,-0.313263), (4733,-0.502257), (4734,-0.211426), (4735,-0.373940), (4736,-0.586159), (4737,-0.252598), (4738,-0.403496), (4739,-0.254342), (4740,-0.418715), (4741,-0.388463), (4742,-0.549124), (4743,-0.292199), (4744,-0.562483), (4745,-0.225202), (4746,-0.377034), (4747,-0.352824), (4748,-0.490254), (4749,-0.598892), (4750,-0.729359), (4751,-0.446887), (4752,-0.605224), (4753,-0.260048), (4754,-0.397947), (4755,-0.256682), (4756,-0.415483), (4757,-0.380121), (4758,-0.541715), (4759,-0.286180), (4760,-0.393886), (4761,-0.443996), (4762,-0.196827), (4763,-0.167972), (4764,-0.326309), (4765,-0.397321), (4766,-0.574700), (4767,-0.291302), (4768,-0.457071), (4769,-0.501139), (4770,-0.279055), (4771,-0.148009), (4772,-0.279872), (4773,-0.320227), (4774,-0.377300), (4775,-0.075323), (4776,-0.435249), (4777,-0.096578), (4778,-0.255379), (4779,-0.236742), (4780,-0.369062), (4781,-0.436361), (4782,-0.606308), (4783,-0.317799), (4784,-0.477527), (4785,-0.158361), (4786,-0.295797), (4787,-0.133167), (4788,-0.293358), (4789,-0.252893), (4790,-0.414017), (4791,-0.152447), (4792,-0.569510), (4793,-0.228980), (4794,-0.430047), (4795,-0.386789), (4796,-0.525152), (4797,-0.630540), (4798,-0.773079), (4799,-0.507332), (4800,-0.663347), (4801,-0.326066), (4802,-0.473721), (4803,-0.353821), (4804,-0.467569), (4805,-0.428494), (4806,-0.555241), (4807,-0.315969), (4808,-0.480812), (4809,-0.142598), (4810,-0.287003), (4811,-0.284159), (4812,-0.451319), (4813,-0.538586), (4814,-0.659767), (4815,-0.422817), (4816,-0.541205), (4817,-0.195102), (4818,-0.370158), (4819,-0.209388), (4820,-0.376084), (4821,-0.338400), (4822,-0.470263), (4823,-0.190577), (4824,-0.410692), (4825,-0.431999), (4826,-0.189946), (4827,-0.221472), (4828,-0.379809), (4829,-0.431773), (4830,-0.586397), (4831,-0.321577), (4832,-0.477128), (4833,-0.532341), (4834,-0.279137), (4835,-0.123006), (4836,-0.306891), (4837,-0.328668), (4838,-0.398283), (4839,-0.136249), (4840,-0.198902), (4841,-0.306144), (4842,0.065970), (4843,-0.112799), (4844,-0.088126), (4845,-0.256683), (4846,-0.335591), (4847,-0.496245), (4848,-0.227248), (4849,-0.379543), (4850,-0.031580), (4851,-0.172265), (4852,-0.022641), (4853,-0.160540), (4854,-0.130288), (4855,-0.308137), (4856,-0.192883), (4857,-0.237884), (4858,-0.010227), (4859,-0.010632), (4860,-0.172219), (4861,-0.213964), (4862,-0.386703), (4863,-0.136285), (4864,-0.262105), (4865,-0.325221), (4866,-0.084089), (4867,0.051597), (4868,-0.093728), (4869,-0.132693), (4870,-0.218101), (4871,0.106174), (4872,-0.146921), (4873,-0.320117), (4874,0.047814), (4875,-0.096121), (4876,-0.082125), (4877,-0.232103), (4878,-0.350954), (4879,-0.501858), (4880,-0.264909), (4881,-0.406064), (4882,-0.124055), (4883,-0.238730), (4884,-0.097002), (4885,-0.260448), (4886,-0.224624), (4887,-0.371815), (4888,-0.403804), (4889,-0.581183), (4890,-0.141719), (4891,-0.294013), (4892,-0.342264), (4893,-0.479237), (4894,-0.218130), (4895,-0.336987), (4896,-0.388024), (4897,-0.540319), (4898,-0.011206), (4899,-0.143996), (4900,-0.193636), (4901,-0.350114), (4902,-0.006797), (4903,-0.119612), (4904,-0.227318), (4905,-0.282538), (4906,-0.049301), (4907,-0.043207), (4908,-0.181106), (4909,-0.277202), (4910,-0.436930), (4911,-0.166536), (4912,-0.341592), (4913,-0.387057), (4914,-0.161723), (4915,-0.023244), (4916,-0.163466), (4917,-0.205674), (4918,-0.255785), (4919,0.035046), (4920,-0.244060), (4921,-0.370344), (4922,0.043110), (4923,-0.105471), (4924,-0.153259), (4925,-0.312060), (4926,-0.080683), (4927,-0.212539), (4928,-0.281228), (4929,-0.424237), (4930,0.116491), (4931,-0.087362), (4932,-0.152801), (4933,-0.295810), (4934,0.062835), (4935,-0.055089), (4936,-0.229218), (4937,-0.315089), (4938,-0.089755), (4939,-0.043711), (4940,-0.228986), (4941,-0.239617), (4942,-0.381229), (4943,-0.124774), (4944,-0.290538), (4945,-0.344831), (4946,-0.134819), (4947,0.002726), (4948,-0.120771), (4949,-0.196893), (4950,-0.257222), (4951,0.015031), (4952,-0.318420), (4953,-0.457246), (4954,-0.052615), (4955,-0.210953), (4956,-0.271276), (4957,-0.421254), (4958,-0.185231), (4959,-0.327313), (4960,-0.395538), (4961,-0.569668), (4962,-0.018250), (4963,-0.187733), (4964,-0.218802), (4965,-0.332081), (4966,0.016809), (4967,-0.154527), (4968,-0.346308), (4969,-0.033649), (4970,-0.178981), (4971,-0.153838), (4972,-0.280592), (4973,-0.383651), (4974,-0.531769), (4975,-0.257656), (4976,-0.402525), (4977,-0.066171), (4978,-0.226832), (4979,-0.086963), (4980,-0.261555), (4981,-0.208542), (4982,-0.378495), (4983,-0.089987), (4984,-0.469887), (4985,-0.156758), (4986,-0.296517), (4987,-0.287167), (4988,-0.457119), (4989,-0.542063), (4990,-0.693895), (4991,-0.431398), (4992,-0.557688), (4993,-0.595719), (4994,-0.346228), (4995,-0.203573), (4996,-0.327070), (4997,-0.354419), (4998,-0.434717), (4999,-0.139240), (5000,-0.413236), (5001,-0.458701), (5002,-0.211069), (5003,-0.235168), (5004,-0.411151), (5005,-0.473340), (5006,-0.622385), (5007,-0.352918), (5008,-0.482922), (5009,-0.563220), (5010,-0.331386), (5011,-0.188261), (5012,-0.343349), (5013,-0.410641), (5014,-0.477934), (5015,-0.194535), (5016,-0.521487), (5017,-0.584133), (5018,-0.293302), (5019,-0.262593), (5020,-0.446471), (5021,-0.482650), (5022,-0.673961), (5023,-0.403104), (5024,-0.608817), (5025,-0.633844), (5026,-0.409436), (5027,-0.221728), (5028,-0.371700), (5029,-0.459431), (5030,-0.496536), (5031,-0.210350), (5032,-0.445331), (5033,-0.222776), (5034,-0.268704), (5035,-0.430761), (5036,-0.395400), (5037,-0.577888), (5038,-0.654936), (5039,-0.803055), (5040,-0.495041), (5041,-0.272024), (5042,-0.337000), (5043,-0.476289), (5044,-0.333170), (5045,-0.382348), (5046,-0.406447), (5047,-0.621446), (5048,-0.356632), (5049,-0.479666), (5050,-0.143776), (5051,-0.315119), (5052,-0.293233), (5053,-0.432058), (5054,-0.516539), (5055,-0.665584), (5056,-0.424921), (5057,-0.551669), (5058,-0.209748), (5059,-0.377372), (5060,-0.240289), (5061,-0.408846), (5062,-0.391136), (5063,-0.539254), (5064,-0.282330), (5065,-0.446240), (5066,-0.077376), (5067,-0.215738), (5068,-0.213820), (5069,-0.360079), (5070,-0.478473), (5071,-0.620085), (5072,-0.350619), (5073,-0.498274), (5074,-0.150311), (5075,-0.311435), (5076,-0.162737), (5077,-0.312715), (5078,-0.273640), (5079,-0.419436), (5080,-0.405909), (5081,-0.544271), (5082,-0.214423), (5083,-0.375547), (5084,-0.350405), (5085,-0.491090), (5086,-0.552347), (5087,-0.721830), (5088,-0.462119), (5089,-0.665515), (5090,-0.299431), (5091,-0.431757), (5092,-0.259372), (5093,-0.431648), (5094,-0.428334), (5095,-0.540685), (5096,-0.287944), (5097,-0.473225), (5098,-0.095532), (5099,-0.255259), (5100,-0.273316), (5101,-0.440482), (5102,-0.495232), (5103,-0.653570), (5104,-0.372494), (5105,-0.540117), (5106,-0.213526), (5107,-0.352352), (5108,-0.197618), (5109,-0.366637), (5110,-0.347068), (5111,-0.477998), (5112,-0.267066), (5113,-0.417970), (5114,-0.067215), (5115,-0.233911), (5116,-0.233860), (5117,-0.366643), (5118,-0.448337), (5119,-0.626186), (5120,-0.299125), (5121,-0.451883), (5122,-0.114139), (5123,-0.245075), (5124,-0.093591), (5125,-0.252392), (5126,-0.171978), (5127,-0.333101), (5128,-0.194159), (5129,-0.368752), (5130,-0.004997), (5131,-0.179126), (5132,-0.159094), (5133,-0.306279), (5134,-0.384260), (5135,-0.545847), (5136,-0.278704), (5137,-0.417066), (5138,-0.122522), (5139,-0.240910), (5140,-0.079676), (5141,-0.273310), (5142,-0.260253), (5143,-0.403725), (5144,-0.189067), (5145,-0.252183), (5146,-0.417953), (5147,0.005263), (5148,-0.144715), (5149,-0.211544), (5150,-0.349907), (5151,-0.092056), (5152,-0.251320), (5153,-0.359958), (5154,-0.516899), (5155,0.059596), (5156,-0.096882), (5157,-0.153028), (5158,-0.279312), (5159,0.073291), (5160,-0.345157), (5161,-0.417565), (5162,-0.175506), (5163,-0.182880), (5164,-0.312420), (5165,-0.364384), (5166,-0.530154), (5167,-0.261151), (5168,-0.398123), (5169,-0.467276), (5170,-0.228930), (5171,-0.070946), (5172,-0.223710), (5173,-0.277534), (5174,-0.349936), (5175,-0.049355), (5176,-0.292695), (5177,-0.351158), (5178,-0.104459), (5179,-0.132735), (5180,-0.291073), (5181,-0.328171), (5182,-0.512520), (5183,-0.217048), (5184,-0.380959), (5185,-0.435709), (5186,-0.210838), (5187,-0.050068), (5188,-0.208869), (5189,-0.260833), (5190,-0.319302), (5191,-0.045196), (5192,-0.332662), (5193,-0.380912), (5194,-0.134670), (5195,-0.149014), (5196,-0.316637), (5197,-0.402051), (5198,-0.579894), (5199,-0.282563), (5200,-0.450186), (5201,-0.529557), (5202,-0.262414), (5203,-0.073773), (5204,-0.244653), (5205,-0.272929), (5206,-0.358806), (5207,-0.077730), (5208,-0.182649), (5209,-0.245295), (5210,-0.421284), (5211,0.005181), (5212,-0.149443), (5213,-0.200944), (5214,-0.371823), (5215,-0.121398), (5216,-0.264870), (5217,-0.284324), (5218,-0.410144), (5219,0.110610), (5220,-0.045868), (5221,-0.112234), (5222,-0.284503), (5223,0.108049), (5224,-0.405162), (5225,-0.063699), (5226,-0.208568), (5227,-0.236844), (5228,-0.334330), (5229,-0.432749), (5230,-0.613841), (5231,-0.318364), (5232,-0.525010), (5233,-0.197022), (5234,-0.328415), (5235,-0.190870), (5236,-0.343164), (5237,-0.325924), (5238,-0.488438), (5239,-0.203180), (5240,-0.360590), (5241,-0.413487), (5242,-0.163532), (5243,-0.142573), (5244,-0.309269), (5245,-0.377488), (5246,-0.563696), (5247,-0.254750), (5248,-0.572873), (5249,-0.637848), (5250,-0.379997), (5251,-0.238269), (5252,-0.378485), (5253,-0.412340), (5254,-0.463841), (5255,-0.225031), (5256,-0.453042), (5257,-0.515695), (5258,-0.267600), (5259,-0.219233), (5260,-0.387326), (5261,-0.475056), (5262,-0.650576), (5263,-0.363000), (5264,-0.515295), (5265,-0.586770), (5266,-0.338212), (5267,-0.182081), (5268,-0.339492), (5269,-0.401675), (5270,-0.494052), (5271,-0.219482), (5272,-0.451669), (5273,-0.613720), (5274,-0.249502), (5275,-0.405979), (5276,-0.377124), (5277,-0.521523), (5278,-0.612509), (5279,-0.795461), (5280,-0.508349), (5281,-0.664827), (5282,-0.305249), (5283,-0.441294), (5284,-0.295383), (5285,-0.448611), (5286,-0.441584), (5287,-0.581806), (5288,-0.345320), (5289,-0.468823), (5290,-0.135719), (5291,-0.298703), (5292,-0.282853), (5293,-0.424465), (5294,-0.512202), (5295,-0.691434), (5296,-0.401073), (5297,-0.551044), (5298,-0.178930), (5299,-0.338658), (5300,-0.181137), (5301,-0.340865), (5302,-0.310156), (5303,-0.487072), (5304,-0.408048), (5305,-0.544550), (5306,-0.219349), (5307,-0.357711), (5308,-0.358123), (5309,-0.512741), (5310,-0.618123), (5311,-0.768564), (5312,-0.488415), (5313,-0.645826), (5314,-0.309472), (5315,-0.446445), (5316,-0.297747), (5317,-0.468626), (5318,-0.420723), (5319,-0.566981), (5320,-0.334678), (5321,-0.492552), (5322,-0.168740), (5323,-0.318249), (5324,-0.318197), (5325,-0.459346), (5326,-0.549863), (5327,-0.718419), (5328,-0.438270), (5329,-0.593821), (5330,-0.256077), (5331,-0.401403), (5332,-0.242493), (5333,-0.376209), (5334,-0.365932), (5335,-0.512190), (5336,-0.485658), (5337,-0.619844), (5338,-0.292319), (5339,-0.445077), (5340,-0.417618), (5341,-0.569913), (5342,-0.637212), (5343,-0.777891), (5344,-0.511217), (5345,-0.645397), (5346,-0.356889), (5347,-0.532414), (5348,-0.372571), (5349,-0.565279), (5350,-0.545715), (5351,-0.682682), (5352,-0.407179), (5353,-0.547401), (5354,-0.192932), (5355,-0.332228), (5356,-0.333566), (5357,-0.487721), (5358,-0.558733), (5359,-0.685480), (5360,-0.441098), (5361,-0.584570), (5362,-0.239857), (5363,-0.409346), (5364,-0.260648), (5365,-0.393901), (5366,-0.342285), (5367,-0.486220), (5368,-0.233478), (5369,-0.383456), (5370,-0.036884), (5371,-0.206836), (5372,-0.225357), (5373,-0.354897), (5374,-0.470961), (5375,-0.589349), (5376,-0.315706), (5377,-0.472184), (5378,-0.120038), (5379,-0.271876), (5380,-0.139897), (5381,-0.293124), (5382,-0.286567), (5383,-0.411924), (5384,-0.304102), (5385,-0.451757), (5386,-0.101008), (5387,-0.248657), (5388,-0.220734), (5389,-0.373956), (5390,-0.424529), (5391,-0.581940), (5392,-0.308760), (5393,-0.467091), (5394,-0.142823), (5395,-0.314159), (5396,-0.166858), (5397,-0.324732), (5398,-0.274048), (5399,-0.423556), (5400,-0.224697), (5401,-0.273874), (5402,-0.457759), (5403,-0.043836), (5404,-0.160833), (5405,-0.225339), (5406,-0.380427), (5407,-0.135581), (5408,-0.305064), (5409,-0.355169), (5410,-0.498641), (5411,0.036509), (5412,-0.089775), (5413,-0.156141), (5414,-0.341416), (5415,0.033954), (5416,-0.401224), (5417,-0.454121), (5418,-0.235286), (5419,-0.220363), (5420,-0.352690), (5421,-0.400477), (5422,-0.555095), (5423,-0.249398), (5424,-0.405412), (5425,-0.449487), (5426,-0.236225), (5427,-0.084741), (5428,-0.221713), (5429,-0.283896), (5430,-0.349335), (5431,-0.070583), (5432,-0.344110), (5433,-0.411872), (5434,-0.179569), (5435,-0.147457), (5436,-0.329952), (5437,-0.379129), (5438,-0.565331), (5439,-0.288438), (5440,-0.429587), (5441,-0.477375), (5442,-0.231602), (5443,-0.068973), (5444,-0.249138), (5445,-0.315504), (5446,-0.400448), (5447,-0.102654), (5448,-0.382217), (5449,-0.427218), (5450,-0.191201), (5451,-0.188357), (5452,-0.338328), (5453,-0.404694), (5454,-0.598335), (5455,-0.318186), (5456,-0.484882), (5457,-0.537316), (5458,-0.323591), (5459,-0.146559), (5460,-0.302574), (5461,-0.374976), (5462,-0.411617), (5463,-0.137041), (5464,-0.226632), (5465,-0.295320), (5466,-0.470383), (5467,-0.056923), (5468,-0.198072), (5469,-0.261651), (5470,-0.439030), (5471,-0.172356), (5472,-0.319541), (5473,-0.370115), (5474,-0.538208), (5475,-0.005376), (5476,-0.149311), (5477,-0.210568), (5478,-0.380514), (5479,0.013898), (5480,-0.369252), (5481,-0.363158), (5482,-0.160585), (5483,-0.088993), (5484,-0.259410), (5485,-0.324379), (5486,-0.503618), (5487,-0.219292), (5488,-0.382269), (5489,-0.456995), (5490,-0.217728), (5491,-0.064848), (5492,-0.208320), (5493,-0.250998), (5494,-0.302968), (5495,-0.029319), (5496,-0.376245), (5497,-0.434245), (5498,-0.172218), (5499,-0.167050), (5500,-0.306803), (5501,-0.362949), (5502,-0.577955), (5503,-0.271795), (5504,-0.496556), (5505,-0.550843), (5506,-0.303681), (5507,-0.146154), (5508,-0.325862), (5509,-0.373180), (5510,-0.446515), (5511,-0.184945), (5512,-0.353501), (5513,-0.495583), (5514,-0.146224), (5515,-0.309671), (5516,-0.260377), (5517,-0.414531), (5518,-0.463246), (5519,-0.605791), (5520,-0.331678), (5521,-0.504881), (5522,-0.178746), (5523,-0.335224), (5524,-0.183746), (5525,-0.349046), (5526,-0.310905), (5527,-0.479924), (5528,-0.404150), (5529,-0.562024), (5530,-0.233566), (5531,-0.365429), (5532,-0.348653), (5533,-0.527891), (5534,-0.601683), (5535,-0.758167), (5536,-0.499846), (5537,-0.609875), (5538,-0.266095), (5539,-0.352899), (5540,-0.255296), (5541,-0.429889), (5542,-0.399644), (5543,-0.536610), (5544,-0.307093), (5545,-0.476112), (5546,-0.168093), (5547,-0.311101), (5548,-0.310580), (5549,-0.448479), (5550,-0.523204), (5551,-0.663427), (5552,-0.386070), (5553,-0.540225), (5554,-0.201085), (5555,-0.343630), (5556,-0.170318), (5557,-0.331905), (5558,-0.312335), (5559,-0.440479), (5560,-0.358675), (5561,-0.528621), (5562,-0.210382), (5563,-0.359897), (5564,-0.356120), (5565,-0.492629), (5566,-0.560385), (5567,-0.712686), (5568,-0.413495), (5569,-0.593197), (5570,-0.222010), (5571,-0.371981), (5572,-0.247441), (5573,-0.415065), (5574,-0.388069), (5575,-0.562661), (5576,-0.304810), (5577,-0.476616), (5578,-0.091497), (5579,-0.242865), (5580,-0.224692), (5581,-0.396035), (5582,-0.465187), (5583,-0.623988), (5584,-0.367990), (5585,-0.513322), (5586,-0.133312), (5587,-0.328806), (5588,-0.176858), (5589,-0.348201), (5590,-0.302157), (5591,-0.428441), (5592,-0.395409), (5593,-0.546314), (5594,-0.221112), (5595,-0.392448), (5596,-0.347338), (5597,-0.507998), (5598,-0.594802), (5599,-0.790296), (5600,-0.502251), (5601,-0.640150), (5602,-0.285682), (5603,-0.472353), (5604,-0.329698), (5605,-0.478743), (5606,-0.445241), (5607,-0.630053), (5608,-0.319716), (5609,-0.493846), (5610,-0.128231), (5611,-0.276813), (5612,-0.282327), (5613,-0.421623), (5614,-0.521896), (5615,-0.668154), (5616,-0.369890), (5617,-0.526368), (5618,-0.165863), (5619,-0.323273), (5620,-0.190368), (5621,-0.310152), (5622,-0.252499), (5623,-0.410836), (5624,-0.177137), (5625,-0.348016), (5626,-0.000053), (5627,-0.173249), (5628,-0.162972), (5629,-0.316200), (5630,-0.393711), (5631,-0.535794), (5632,-0.307203), (5633,-0.461827), (5634,-0.108285), (5635,-0.267549), (5636,-0.116998), (5637,-0.285091), (5638,-0.258089), (5639,-0.362081), (5640,-0.238931), (5641,-0.382403), (5642,-0.060452), (5643,-0.220185), (5644,-0.228950), (5645,-0.404939), (5646,-0.450867), (5647,-0.599448), (5648,-0.342993), (5649,-0.514800), (5650,-0.171013), (5651,-0.308912), (5652,-0.161148), (5653,-0.334814), (5654,-0.294343), (5655,-0.443851), (5656,-0.243601), (5657,-0.309967), (5658,-0.439970), (5659,-0.059027), (5660,-0.189494), (5661,-0.266078), (5662,-0.391436), (5663,-0.137298), (5664,-0.297025), (5665,-0.360604), (5666,-0.511509), (5667,0.047798), (5668,-0.142587), (5669,-0.175972), (5670,-0.329663), (5671,0.028982), (5672,-0.339773), (5673,-0.409388), (5674,-0.149677), (5675,-0.147766), (5676,-0.321425), (5677,-0.387328), (5678,-0.606980), (5679,-0.298497), (5680,-0.454974), (5681,-0.522273), (5682,-0.274171), (5683,-0.120370), (5684,-0.267556), (5685,-0.359469), (5686,-0.433267), (5687,-0.141973), (5688,-0.425719), (5689,-0.491621), (5690,-0.239343), (5691,-0.182153), (5692,-0.317730), (5693,-0.380846), (5694,-0.546615), (5695,-0.262753), (5696,-0.416445), (5697,-0.488847), (5698,-0.212417), (5699,-0.063256), (5700,-0.258750), (5701,-0.301428), (5702,-0.351539), (5703,-0.061171), (5704,-0.321698), (5705,-0.354621), (5706,-0.114885), (5707,-0.143161), (5708,-0.300101), (5709,-0.356248), (5710,-0.517372), (5711,-0.261381), (5712,-0.406706), (5713,-0.487010), (5714,-0.270035), (5715,-0.093930), (5716,-0.222544), (5717,-0.254533), (5718,-0.331118), (5719,-0.076516), (5720,-0.176795), (5721,-0.224113), (5722,-0.369908), (5723,0.028217), (5724,-0.136620), (5725,-0.157000), (5726,-0.334379), (5727,-0.077925), (5728,-0.213964), (5729,-0.264538), (5730,-0.433088), (5731,0.115537), (5732,-0.040014), (5733,-0.107777), (5734,-0.269827), (5735,0.130158), (5736,-0.218152), (5737,-0.287304), (5738,-0.052678), (5739,-0.042871), (5740,-0.200275), (5741,-0.232734), (5742,-0.404540), (5743,-0.112318), (5744,-0.262753), (5745,-0.336552), (5746,-0.099602), (5747,0.045839), (5748,-0.104139), (5749,-0.172358), (5750,-0.262881), (5751,0.029347), (5752,-0.296209), (5753,-0.365361), (5754,-0.104260), (5755,-0.112561), (5756,-0.257893), (5757,-0.314967), (5758,-0.511857), (5759,-0.227532), (5760,-0.425812), (5761,-0.590186), (5762,-0.238510), (5763,-0.401487), (5764,-0.242113), (5765,-0.387438), (5766,-0.368339), (5767,-0.527139), (5768,-0.341285), (5769,-0.526560), (5770,-0.190676), (5771,-0.332288), (5772,-0.281141), (5773,-0.419034), (5774,-0.507698), (5775,-0.661389), (5776,-0.371491), (5777,-0.522389), (5778,-0.180469), (5779,-0.332763), (5780,-0.219832), (5781,-0.348909), (5782,-0.351637), (5783,-0.486287), (5784,-0.429097), (5785,-0.581392), (5786,-0.248294), (5787,-0.413131), (5788,-0.410750), (5789,-0.571410), (5790,-0.625697), (5791,-0.769639), (5792,-0.474625), (5793,-0.607415), (5794,-0.289646), (5795,-0.431721), (5796,-0.274664), (5797,-0.485487), (5798,-0.432017), (5799,-0.577812), (5800,-0.340862), (5801,-0.498730), (5802,-0.156810), (5803,-0.303532), (5804,-0.317412), (5805,-0.455305), (5806,-0.519817), (5807,-0.663753), (5808,-0.400792), (5809,-0.523363), (5810,-0.206520), (5811,-0.383436), (5812,-0.247744), (5813,-0.394472), (5814,-0.353538), (5815,-0.489114), (5816,-0.395694), (5817,-0.563318), (5818,-0.200953), (5819,-0.358364), (5820,-0.362952), (5821,-0.518496), (5822,-0.584399), (5823,-0.749242), (5824,-0.521578), (5825,-0.676202), (5826,-0.277144), (5827,-0.437335), (5828,-0.283997), (5829,-0.453481), (5830,-0.430198), (5831,-0.549982), (5832,-0.286095), (5833,-0.448145), (5834,-0.112725), (5835,-0.273842), (5836,-0.264961), (5837,-0.424225), (5838,-0.498024), (5839,-0.657288), (5840,-0.370176), (5841,-0.517831), (5842,-0.194019), (5843,-0.358856), (5844,-0.199476), (5845,-0.324833), (5846,-0.281582), (5847,-0.458961), (5848,-0.472372), (5849,-0.638605), (5850,-0.290642), (5851,-0.409030), (5852,-0.440099), (5853,-0.592857), (5854,-0.685234), (5855,-0.809664), (5856,-0.508150), (5857,-0.658128), (5858,-0.287404), (5859,-0.448991), (5860,-0.355102), (5861,-0.481855), (5862,-0.440458), (5863,-0.607618), (5864,-0.639613), (5865,-0.375256), (5866,-0.115082), (5867,-0.199563), (5868,-0.356510), (5869,-0.331368), (5870,-0.486919), (5871,-0.528200), (5872,-0.699080), (5873,-0.436119), (5874,-0.205206), (5875,-0.298515), (5876,-0.426195), (5877,-0.264492), (5878,-0.339681), (5879,-0.379109), (5880,-0.124044), (5881,-0.289345), (5882,-0.337132), (5883,-0.094146), (5884,-0.096411), (5885,-0.252425), (5886,-0.303463), (5887,-0.484561), (5888,-0.230423), (5889,-0.409662), (5890,-0.434688), (5891,-0.201452), (5892,-0.040682), (5893,-0.199019), (5894,-0.259348), (5895,-0.315495), (5896,-0.491478), (5897,-0.232237), (5898,-0.368739), (5899,-0.037495), (5900,-0.176327), (5901,-0.203207), (5902,-0.337393), (5903,-0.398649), (5904,-0.543975), (5905,-0.248040), (5906,-0.427273), (5907,-0.100218), (5908,-0.253439), (5909,-0.079664), (5910,-0.228245), (5911,-0.208212), (5912,-0.220696), (5913,-0.304714), (5914,-0.491385), (5915,-0.046341), (5916,-0.212111), (5917,-0.258039), (5918,-0.434955), (5919,-0.190572), (5920,-0.312216), (5921,-0.376722), (5922,-0.553175), (5923,-0.016629), (5924,-0.170314), (5925,-0.219961), (5926,-0.338812), (5927,0.009151), (5928,-0.290394), (5929,-0.476132), (5930,-0.138858), (5931,-0.280470), (5932,-0.257651), (5933,-0.400660), (5934,-0.484677), (5935,-0.633722), (5936,-0.369835), (5937,-0.532348), (5938,-0.172307), (5939,-0.346436), (5940,-0.190775), (5941,-0.355612), (5942,-0.314215), (5943,-0.470229), (5944,-0.247681), (5945,-0.322870), (5946,-0.487243), (5947,-0.062174), (5948,-0.220975), (5949,-0.265049), (5950,-0.402479), (5951,-0.155780), (5952,-0.323866), (5953,-0.417639), (5954,-0.570404), (5955,-0.063119), (5956,-0.205195), (5957,-0.244623), (5958,-0.382985), (5959,-0.005755), (5960,-0.160843), (5961,-0.314064), (5962,-0.360925), (5963,-0.087745), (5964,-0.075145), (5965,-0.239055), (5966,-0.271977), (5967,-0.463758), (5968,-0.207767), (5969,-0.338234), (5970,-0.451975), (5971,-0.201557), (5972,-0.033817), (5973,-0.213983), (5974,-0.254338), (5975,-0.359720), (5976,-0.258868), (5977,-0.322910), (5978,-0.462206), (5979,-0.075220), (5980,-0.213120), (5981,-0.270199), (5982,-0.411348), (5983,-0.145138), (5984,-0.322054), (5985,-0.360549), (5986,-0.469181), (5987,0.074798), (5988,-0.077961), (5989,-0.125285), (5990,-0.309170), (5991,0.027184), (5992,-0.214296), (5993,-0.385175), (5994,-0.056724), (5995,-0.199726), (5996,-0.174127), (5997,-0.315739), (5998,-0.403933), (5999,-0.549728), (6000,-0.284914), (6001,-0.420484), (6002,-0.066948), (6003,-0.225285), (6004,-0.048723), (6005,-0.261399), (6006,-0.225581), (6007,-0.385308), (6008,-0.303504), (6009,-0.447440), (6010,-0.073466), (6011,-0.242479), (6012,-0.226629), (6013,-0.400295), (6014,-0.441577), (6015,-0.588768), (6016,-0.634696), (6017,-0.706171), (6018,-0.458076), (6019,-0.310311), (6020,-0.465392), (6021,-0.536868), (6022,-0.600910), (6023,-0.292427), (6024,-0.476312), (6025,-0.639759), (6026,-0.274608), (6027,-0.415294), (6028,-0.404553), (6029,-0.576359), (6030,-0.656664), (6031,-0.808958), (6032,-0.507908), (6033,-0.669958), (6034,-0.330361), (6035,-0.471510), (6036,-0.329782), (6037,-0.492295), (6038,-0.467159), (6039,-0.618991), (6040,-0.357420), (6041,-0.505075), (6042,-0.543570), (6043,-0.296871), (6044,-0.275442), (6045,-0.438426), (6046,-0.485750), (6047,-0.661269), (6048,-0.397382), (6049,-0.534811), (6050,-0.598854), (6051,-0.324747), (6052,-0.186269), (6053,-0.354362), (6054,-0.407259), (6055,-0.473161), (6056,-0.350938), (6057,-0.527854), (6058,-0.168282), (6059,-0.281097), (6060,-0.328884), (6061,-0.498830), (6062,-0.598640), (6063,-0.772769), (6064,-0.462426), (6065,-0.629593), (6066,-0.289989), (6067,-0.430675), (6068,-0.267112), (6069,-0.418949), (6070,-0.405886), (6071,-0.560040), (6072,-0.530722), (6073,-0.670011), (6074,-0.313689), (6075,-0.458087), (6076,-0.438524), (6077,-0.611721), (6078,-0.695738), (6079,-0.846179), (6080,-0.567427), (6081,-0.736446), (6082,-0.365722), (6083,-0.542638), (6084,-0.398123), (6085,-0.561100), (6086,-0.524349), (6087,-0.643670), (6088,-0.415079), (6089,-0.549265), (6090,-0.238459), (6091,-0.372176), (6092,-0.394879), (6093,-0.539284), (6094,-0.626551), (6095,-0.747725), (6096,-0.475473), (6097,-0.614768), (6098,-0.275165), (6099,-0.445581), (6100,-0.309425), (6101,-0.453361), (6102,-0.431474), (6103,-0.600024), (6104,-0.315699), (6105,-0.485182), (6106,-0.525537), (6107,-0.284411), (6108,-0.281103), (6109,-0.458482), (6110,-0.522988), (6111,-0.701763), (6112,-0.444376), (6113,-0.579019), (6114,-0.632849), (6115,-0.401009), (6116,-0.284364), (6117,-0.417148), (6118,-0.465399), (6119,-0.522942), (6120,-0.213532), (6121,-0.363973), (6122,-0.386676), (6123,-0.142758), (6124,-0.139913), (6125,-0.306146), (6126,-0.362293), (6127,-0.541532), (6128,-0.241408), (6129,-0.379771), (6130,-0.443820), (6131,-0.199901), (6132,-0.030302), (6133,-0.183993), (6134,-0.243396), (6135,-0.332516), (6136,-0.089994), (6137,-0.247404), (6138,-0.304015), (6139,-0.098649), (6140,-0.062361), (6141,-0.231380), (6142,-0.301929), (6143,-0.496033), (6144,-0.651114), (6145,-0.364466), (6146,-0.554850), (6147,-0.217106), (6148,-0.364298), (6149,-0.224893), (6150,-0.354889), (6151,-0.335326), (6152,-0.625578), (6153,-0.367727), (6154,-0.522808), (6155,-0.171596), (6156,-0.356871), (6157,-0.364715), (6158,-0.509577), (6159,-0.551792), (6160,-0.726384), (6161,-0.450881), (6162,-0.589244), (6163,-0.297023), (6164,-0.446067), (6165,-0.279718), (6166,-0.429696), (6167,-0.409200), (6168,-0.407289), (6169,-0.575839), (6170,-0.645924), (6171,-0.415010), (6172,-0.412166), (6173,-0.585368), (6174,-0.606212), (6175,-0.790560), (6176,-0.520167), (6177,-0.657603), (6178,-0.711426), (6179,-0.479586), (6180,-0.347150), (6181,-0.508274), (6182,-0.546769), (6183,-0.605702), (6184,-0.336236), (6185,-0.500146), (6186,-0.567445), (6187,-0.333282), (6188,-0.290957), (6189,-0.432570), (6190,-0.479894), (6191,-0.682357), (6192,-0.368764), (6193,-0.550790), (6194,-0.587888), (6195,-0.341189), (6196,-0.192492), (6197,-0.355012), (6198,-0.417658), (6199,-0.497493), (6200,-0.316748), (6201,-0.476945), (6202,-0.527982), (6203,-0.269204), (6204,-0.273793), (6205,-0.438166), (6206,-0.485947), (6207,-0.656363), (6208,-0.410591), (6209,-0.578214), (6210,-0.634361), (6211,-0.375583), (6212,-0.211094), (6213,-0.369894), (6214,-0.445546), (6215,-0.494267), (6216,-0.288437), (6217,-0.447701), (6218,-0.499202), (6219,-0.280367), (6220,-0.266840), (6221,-0.402417), (6222,-0.481788), (6223,-0.656380), (6224,-0.346044), (6225,-0.501595), (6226,-0.566564), (6227,-0.309177), (6228,-0.162808), (6229,-0.305811), (6230,-0.363817), (6231,-0.426933), (6232,-0.310752), (6233,-0.474663), (6234,-0.535919), (6235,-0.303152), (6236,-0.291479), (6237,-0.445170), (6238,-0.524541), (6239,-0.681952), (6240,-0.411558), (6241,-0.563390), (6242,-0.618146), (6243,-0.401172), (6244,-0.245968), (6245,-0.376904), (6246,-0.452556), (6247,-0.544933), (6248,-0.487743), (6249,-0.627039), (6250,-0.255382), (6251,-0.444376), (6252,-0.430849), (6253,-0.563176), (6254,-0.660199), (6255,-0.809244), (6256,-0.520735), (6257,-0.662811), (6258,-0.326927), (6259,-0.490837), (6260,-0.319378), (6261,-0.487008), (6262,-0.473944), (6263,-0.628099), (6264,-0.343310), (6265,-0.505824), (6266,-0.543392), (6267,-0.312016), (6268,-0.249717), (6269,-0.419663), (6270,-0.483242), (6271,-0.677810), (6272,-0.596005), (6273,-0.744117), (6274,-0.366894), (6275,-0.519658), (6276,-0.394185), (6277,-0.541840), (6278,-0.511588), (6279,-0.662956), (6280,-0.472919), (6281,-0.652627), (6282,-0.333462), (6283,-0.461142), (6284,-0.442036), (6285,-0.590154), (6286,-0.673245), (6287,-0.793956), (6288,-0.539355), (6289,-0.724629), (6290,-0.357162), (6291,-0.489482), (6292,-0.382593), (6293,-0.525139), (6294,-0.496283), (6295,-0.643468), (6296,-0.827353), (6297,-0.562533), (6298,-0.320937), (6299,-0.345963), (6300,-0.535421), (6301,-0.493560), (6302,-0.654220), (6303,-0.712227), (6304,-0.874741), (6305,-0.569977), (6306,-0.354392), (6307,-0.409149), (6308,-0.549365), (6309,-0.416929), (6310,-0.472149), (6311,-0.597506), (6312,-1.000631), (6313,-0.315439), (6314,-0.467277), (6315,-0.527600), (6316,-0.667823), (6317,-0.689599), (6318,-0.816809), (6319,-0.885498), (6320,-1.039659), (6321,-0.377692), (6322,-0.527670), (6323,-0.556873), (6324,-0.693382), (6325,-0.459219), (6326,-0.598971), (6327,-0.678812), (6328,-0.871520), (6329,-0.569543), (6330,-0.302399), (6331,-0.377588), (6332,-0.518743), (6333,-0.517752), (6334,-0.712319), (6335,-0.761967), (6336,-0.902652), (6337,-0.631326), (6338,-0.412028), (6339,-0.449596), (6340,-0.614440), (6341,-0.488966), (6342,-0.535358), (6343,-0.551561), (6344,-0.739159), (6345,-0.468766), (6346,-0.235066), (6347,-0.274958), (6348,-0.478348), (6349,-0.470394), (6350,-0.663107), (6351,-0.707175), (6352,-0.850647), (6353,-0.582577), (6354,-0.332622), (6355,-0.366008), (6356,-0.528528), (6357,-0.381227), (6358,-0.446196), (6359,-0.503269), (6360,-0.808850), (6361,-0.520811), (6362,-0.254595), (6363,-0.354404), (6364,-0.513205), (6365,-0.468094), (6366,-0.647333), (6367,-0.665853), (6368,-0.868780), (6369,-0.573309), (6370,-0.345182), (6371,-0.451497), (6372,-0.602402), (6373,-0.455100), (6374,-0.520070), (6375,-0.542310), (6376,-0.678349), (6377,-0.411212), (6378,-0.191444), (6379,-0.270816), (6380,-0.418470), (6381,-0.397048), (6382,-0.581396), (6383,-0.627787), (6384,-0.765223), (6385,-0.512944), (6386,-0.277385), (6387,-0.321459), (6388,-0.469577), (6389,-0.320880), (6390,-0.399788), (6391,-0.450362), (6392,-0.718779), (6393,-0.431667), (6394,-0.195181), (6395,-0.263870), (6396,-0.433353), (6397,-0.386846), (6398,-0.580486), (6399,-0.659394), (6400,-0.804256), (6401,-0.522717), (6402,-0.270439), (6403,-0.330769), (6404,-0.488173), (6405,-0.346445), (6406,-0.417457), (6407,-0.493578), (6408,-0.820060), (6409,-0.523656), (6410,-0.279274), (6411,-0.350749), (6412,-0.503977), (6413,-0.489523), (6414,-0.690590), (6415,-0.741627), (6416,-0.903678), (6417,-0.612383), (6418,-0.375903), (6419,-0.408362), (6420,-0.556943), (6421,-0.425434), (6422,-0.528493), (6423,-0.575817), (6424,-0.370915), (6425,-0.499992), (6426,-0.575643), (6427,-0.302000), (6428,-0.295443), (6429,-0.466779), (6430,-0.518286), (6431,-0.704024), (6432,-0.420162), (6433,-0.581286), (6434,-0.609099), (6435,-0.371222), (6436,-0.228098), (6437,-0.403154), (6438,-0.437009), (6439,-0.539141), (6440,-0.410418), (6441,-0.565036), (6442,-0.215214), (6443,-0.355899), (6444,-0.353524), (6445,-0.482595), (6446,-0.602379), (6447,-0.741668), (6448,-0.464312), (6449,-0.621716), (6450,-0.300228), (6451,-0.434414), (6452,-0.268064), (6453,-0.446840), (6454,-0.422630), (6455,-0.569352), (6456,-0.483365), (6457,-0.647276), (6458,-0.299776), (6459,-0.454394), (6460,-0.426002), (6461,-0.607100), (6462,-0.698087), (6463,-0.857351), (6464,-0.595317), (6465,-0.726710), (6466,-0.380144), (6467,-0.520829), (6468,-0.398143), (6469,-0.545334), (6470,-0.533198), (6471,-0.647872), (6472,-0.491748), (6473,-0.621282), (6474,-0.294220), (6475,-0.432120), (6476,-0.395832), (6477,-0.589935), (6478,-0.646082), (6479,-0.820675), (6480,-0.523344), (6481,-0.676102), (6482,-0.310024), (6483,-0.473934), (6484,-0.367509), (6485,-0.504012), (6486,-0.458901), (6487,-0.614915), (6488,-0.320834), (6489,-0.465233), (6490,-0.545531), (6491,-0.273284), (6492,-0.286695), (6493,-0.452929), (6494,-0.519758), (6495,-0.671589), (6496,-0.372398), (6497,-0.551174), (6498,-0.609644), (6499,-0.355975), (6500,-0.180803), (6501,-0.343780), (6502,-0.392964), (6503,-0.485341), (6504,-0.561926), (6505,-0.314294), (6506,-0.381123), (6507,-0.527382), (6508,-0.507818), (6509,-0.700989), (6510,-0.755276), (6511,-0.934979), (6512,-0.630215), (6513,-0.371901), (6514,-0.431297), (6515,-0.565013), (6516,-0.400994), (6517,-0.460390), (6518,-0.557413), (6519,-0.702745), (6520,-0.410054), (6521,-0.586969), (6522,-0.238080), (6523,-0.395948), (6524,-0.411224), (6525,-0.546794), (6526,-0.668901), (6527,-0.798905), (6528,-0.619086), (6529,-0.775564), (6530,-0.455009), (6531,-0.621242), (6532,-0.452569), (6533,-0.579786), (6534,-0.546285), (6535,-0.716701), (6536,-0.523414), (6537,-0.680355), (6538,-0.320776), (6539,-0.486546), (6540,-0.497640), (6541,-0.640179), (6542,-0.711655), (6543,-0.838408), (6544,-0.572191), (6545,-0.740284), (6546,-0.413686), (6547,-0.576206), (6548,-0.427972), (6549,-0.564481), (6550,-0.545375), (6551,-0.686994), (6552,-0.849044), (6553,-0.580974), (6554,-0.337518), (6555,-0.406207), (6556,-0.538070), (6557,-0.513861), (6558,-0.722361), (6559,-0.760856), (6560,-0.907577), (6561,-0.631611), (6562,-0.402094), (6563,-0.433626), (6564,-0.613329), (6565,-0.479960), (6566,-0.558404), (6567,-0.623374), (6568,-1.039504), (6569,-0.349209), (6570,-0.497327), (6571,-0.545115), (6572,-0.701129), (6573,-0.716400), (6574,-0.886346), (6575,-0.929487), (6576,-1.095257), (6577,-0.412858), (6578,-0.577232), (6579,-0.650567), (6580,-0.805648), (6581,-0.570558), (6582,-0.691269), (6583,-0.742306), (6584,-0.940123), (6585,-0.660907), (6586,-0.397483), (6587,-0.438765), (6588,-0.584097), (6589,-0.619342), (6590,-0.804617), (6591,-0.870983), (6592,-1.007022), (6593,-0.744525), (6594,-0.499216), (6595,-0.546070), (6596,-0.696975), (6597,-0.516694), (6598,-0.577487), (6599,-0.622951), (6600,-0.824951), (6601,-0.561527), (6602,-0.314358), (6603,-0.383047), (6604,-0.555780), (6605,-0.527851), (6606,-0.695017), (6607,-0.737226), (6608,-0.873735), (6609,-0.615414), (6610,-0.351990), (6611,-0.426715), (6612,-0.578553), (6613,-0.434038), (6614,-0.530591), (6615,-0.566770), (6616,-0.890929), (6617,-0.578732), (6618,-0.365007), (6619,-0.402112), (6620,-0.553944), (6621,-0.517192), (6622,-0.712223), (6623,-0.768370), (6624,-0.924847), (6625,-0.632626), (6626,-0.391030), (6627,-0.463432), (6628,-0.641744), (6629,-0.470285), (6630,-0.551980), (6631,-0.626711), (6632,-0.794798), (6633,-0.499790), (6634,-0.263304), (6635,-0.316201), (6636,-0.491720), (6637,-0.452182), (6638,-0.642103), (6639,-0.701500), (6640,-0.858910), (6641,-0.563433), (6642,-0.326483), (6643,-0.361729), (6644,-0.522852), (6645,-0.389483), (6646,-0.446100), (6647,-0.502246), (6648,-0.777633), (6649,-0.506313), (6650,-0.288869), (6651,-0.342229), (6652,-0.444825), (6653,-0.439194), (6654,-0.616579), (6655,-0.668543), (6656,-0.824557), (6657,-0.514215), (6658,-0.270302), (6659,-0.331558), (6660,-0.510797), (6661,-0.375105), (6662,-0.448903), (6663,-0.509233), (6664,-0.831069), (6665,-0.507257), (6666,-0.309794), (6667,-0.362227), (6668,-0.516382), (6669,-0.512141), (6670,-0.679301), (6671,-0.737307), (6672,-0.908187), (6673,-0.580199), (6674,-0.358108), (6675,-0.449095), (6676,-0.582348), (6677,-0.431333), (6678,-0.521387), (6679,-0.559882), (6680,-0.350803), (6681,-0.537011), (6682,-0.601054), (6683,-0.347843), (6684,-0.275324), (6685,-0.448527), (6686,-0.539977), (6687,-0.711783), (6688,-0.419555), (6689,-0.565351), (6690,-0.617784), (6691,-0.362256), (6692,-0.209382), (6693,-0.369109), (6694,-0.395526), (6695,-0.503231), (6696,-0.374978), (6697,-0.557466), (6698,-0.218790), (6699,-0.368304), (6700,-0.357100), (6701,-0.510322), (6702,-0.575298), (6703,-0.719696), (6704,-0.462778), (6705,-0.619256), (6706,-0.284762), (6707,-0.432880), (6708,-0.278146), (6709,-0.442520), (6710,-0.417841), (6711,-0.574325), (6712,-0.503660), (6713,-0.636913), (6714,-0.315894), (6715,-0.452860), (6716,-0.476027), (6717,-0.613463), (6718,-0.698870), (6719,-0.855817), (6720,-0.590997), (6721,-0.783241), (6722,-0.411121), (6723,-0.596402), (6724,-0.464429), (6725,-0.624157), (6726,-0.534914), (6727,-0.662594), (6728,-0.525048), (6729,-0.675490), (6730,-0.340069), (6731,-0.484931), (6732,-0.498812), (6733,-0.660862), (6734,-0.751379), (6735,-0.891138), (6736,-0.619818), (6737,-0.741919), (6738,-0.425546), (6739,-0.553690), (6740,-0.369689), (6741,-0.525703), (6742,-0.507993), (6743,-0.681196), (6744,-0.339739), (6745,-0.511545), (6746,-0.581624), (6747,-0.323773), (6748,-0.334861), (6749,-0.492734), (6750,-0.514974), (6751,-0.686780), (6752,-0.391303), (6753,-0.558469), (6754,-0.598818), (6755,-0.350259), (6756,-0.189026), (6757,-0.361758), (6758,-0.409546), (6759,-0.481484), (6760,-0.544600), (6761,-0.293712), (6762,-0.380053), (6763,-0.501697), (6764,-0.502102), (6765,-0.656257), (6766,-0.688252), (6767,-0.871204), (6768,-0.594774), (6769,-0.384299), (6770,-0.413972), (6771,-0.585778), (6772,-0.441726), (6773,-0.514135), (6774,-0.588396), (6775,-0.748587), (6776,-0.511637), (6777,-0.647214), (6778,-0.319225), (6779,-0.457588), (6780,-0.464499), (6781,-0.608898), (6782,-0.681306), (6783,-0.853576), (6784,-1.145218), (6785,-0.424266), (6786,-0.587249), (6787,-0.662438), (6788,-0.809166), (6789,-0.568960), (6790,-0.738450), (6791,-0.782054), (6792,-1.037003), (6793,-0.367610), (6794,-0.532910), (6795,-0.609964), (6796,-0.734852), (6797,-0.734800), (6798,-0.907069), (6799,-0.927913), (6800,-1.090433), (6801,-0.452160), (6802,-0.606315), (6803,-0.622975), (6804,-0.815689), (6805,-0.569911), (6806,-0.688298), (6807,-0.752811), (6808,-0.894423), (6809,-0.623103), (6810,-0.379648), (6811,-0.425112), (6812,-0.586236), (6813,-0.555990), (6814,-0.767276), (6815,-0.815527), (6816,-0.952030), (6817,-0.695575), (6818,-0.455839), (6819,-0.545429), (6820,-0.684255), (6821,-0.547636), (6822,-0.617722), (6823,-0.644601), (6824,-0.870752), (6825,-0.566452), (6826,-0.267262), (6827,-0.436281), (6828,-0.501720), (6829,-0.684672), (6830,-0.674858), (6831,-0.813221), (6832,-0.867514), (6833,-0.608267), (6834,-0.362031), (6835,-0.530118), (6836,-0.574655), (6837,-0.639625), (6838,-0.474672), (6839,-0.645551), (6840,-1.066791), (6841,-0.408080), (6842,-0.560381), (6843,-0.619315), (6844,-0.785078), (6845,-0.790599), (6846,-0.954973), (6847,-0.986968), (6848,-1.143446), (6849,-0.459187), (6850,-0.602659), (6851,-0.672275), (6852,-0.855697), (6853,-0.627570), (6854,-0.774291), (6855,-0.855059), (6856,-0.947899), (6857,-0.698877), (6858,-0.426624), (6859,-0.602150), (6860,-0.656437), (6861,-0.796659), (6862,-0.820289), (6863,-0.942860), (6864,-0.993433), (6865,-0.749051), (6866,-0.488414), (6867,-0.627240), (6868,-0.686173), (6869,-0.752539), (6870,-0.586659), (6871,-0.748709), (6872,-0.951636), (6873,-0.667311), (6874,-0.403423), (6875,-0.455851), (6876,-0.621157), (6877,-0.579296), (6878,-0.791045), (6879,-0.858338), (6880,-1.026431), (6881,-0.740709), (6882,-0.526057), (6883,-0.556193), (6884,-0.697342), (6885,-0.537962), (6886,-0.626162), (6887,-0.685096), (6888,-0.733810), (6889,-0.868922), (6890,-0.194883), (6891,-0.351361), (6892,-0.404257), (6893,-0.561198), (6894,-0.580188), (6895,-0.751525), (6896,-0.834152), (6897,-0.981337), (6898,-0.290579), (6899,-0.434515), (6900,-0.485089), (6901,-0.647602), (6902,-0.412049), (6903,-0.541589), (6904,-0.751479), (6905,-0.469940), (6906,-0.232063), (6907,-0.266845), (6908,-0.437255), (6909,-0.404217), (6910,-0.602967), (6911,-0.650291), (6912,-0.834169), (6913,-0.543808), (6914,-0.301749), (6915,-0.334208), (6916,-0.516696), (6917,-0.354530), (6918,-0.441797), (6919,-0.473792), (6920,-0.709699), (6921,-0.874073), (6922,-0.179132), (6923,-0.336073), (6924,-0.399652), (6925,-0.539874), (6926,-0.535170), (6927,-0.704653), (6928,-0.751044), (6929,-0.877798), (6930,-0.215374), (6931,-0.352340), (6932,-0.416846), (6933,-0.589585), (6934,-0.356348), (6935,-0.464524), (6936,-0.833735), (6937,-0.576347), (6938,-0.332435), (6939,-0.395081), (6940,-0.571533), (6941,-0.531532), (6942,-0.744678), (6943,-0.808257), (6944,-0.959625), (6945,-0.679940), (6946,-0.466221), (6947,-0.524221), (6948,-0.669090), (6949,-0.475803), (6950,-0.533346), (6951,-0.600638), (6952,-0.789633), (6953,-0.549427), (6954,-0.289259), (6955,-0.341223), (6956,-0.487481), (6957,-0.461412), (6958,-0.634145), (6959,-0.696798), (6960,-0.845380), (6961,-0.570340), (6962,-0.329677), (6963,-0.384897), (6964,-0.530693), (6965,-0.365740), (6966,-0.434892), (6967,-0.508690), (6968,-0.771535), (6969,-0.488136), (6970,-0.251187), (6971,-0.315229), (6972,-0.494931), (6973,-0.465613), (6974,-0.653680), (6975,-0.710754), (6976,-0.882560), (6977,-0.590338), (6978,-0.321335), (6979,-0.360300), (6980,-0.512131), (6981,-0.372726), (6982,-0.471602), (6983,-0.519390), (6984,-0.810575), (6985,-0.533212), (6986,-0.292086), (6987,-0.345447), (6988,-0.472194), (6989,-0.462850), (6990,-0.662057), (6991,-0.706594), (6992,-0.851926), (6993,-0.555985), (6994,-0.324145), (6995,-0.361244), (6996,-0.532123), (6997,-0.378786), (6998,-0.437719), (6999,-0.492469), (7000,-0.841249), (7001,-0.577362), (7002,-0.311615), (7003,-0.358006), (7004,-0.521453), (7005,-0.526504), (7006,-0.682518), (7007,-0.719154), (7008,-0.873308), (7009,-0.581087), (7010,-0.354356), (7011,-0.417472), (7012,-0.618539), (7013,-0.452660), (7014,-0.500910), (7015,-0.549161), (7016,-0.817579), (7017,-0.181166), (7018,-0.319991), (7019,-0.372425), (7020,-0.511714), (7021,-0.531168), (7022,-0.689042), (7023,-0.735433), (7024,-0.936500), (7025,-0.252711), (7026,-0.397109), (7027,-0.449543), (7028,-0.612520), (7029,-0.378827), (7030,-0.506970), (7031,-0.545929), (7032,-0.942084), (7033,-0.272228), (7034,-0.444960), (7035,-0.483462), (7036,-0.640403), (7037,-0.662642), (7038,-0.832126), (7039,-0.875730), (7040,-1.075870), (7041,-0.831488), (7042,-0.610800), (7043,-0.625138), (7044,-0.790444), (7045,-0.630137), (7046,-0.686747), (7047,-0.748004), (7048,-0.894726), (7049,-1.009864), (7050,-0.344190), (7051,-0.502990), (7052,-0.564710), (7053,-0.703073), (7054,-0.716020), (7055,-0.861352), (7056,-0.896597), (7057,-1.077226), (7058,-0.385071), (7059,-0.572676), (7060,-0.619067), (7061,-0.761606), (7062,-0.528376), (7063,-0.676957), (7064,-0.954204), (7065,-1.121827), (7066,-0.435252), (7067,-0.608911), (7068,-0.659022), (7069,-0.781129), (7070,-0.779675), (7071,-0.948694), (7072,-1.040608), (7073,-1.186866), (7074,-0.529088), (7075,-0.644226), (7076,-0.704550), (7077,-0.871716), (7078,-0.602713), (7079,-0.769879), (7080,-0.874328), (7081,-1.017337), (7082,-0.358626), (7083,-0.487703), (7084,-0.552672), (7085,-0.725875), (7086,-0.740682), (7087,-0.869752), (7088,-0.930081), (7089,-1.081449), (7090,-0.393008), (7091,-0.549955), (7092,-0.628863), (7093,-0.810419), (7094,-0.602736), (7095,-0.739702), (7096,-1.009053), (7097,-1.159494), (7098,-0.473376), (7099,-0.607099), (7100,-0.670208), (7101,-0.811357), (7102,-0.845676), (7103,-0.960814), (7104,-1.009065), (7105,-1.169255), (7106,-0.507295), (7107,-0.608500), (7108,-0.681366), (7109,-0.819728), (7110,-0.582785), (7111,-0.767597), (7112,-0.839535), (7113,-0.980684), (7114,-0.321973), (7115,-0.458940), (7116,-0.525305), (7117,-0.677606), (7118,-0.661757), (7119,-0.795010), (7120,-0.864625), (7121,-1.030858), (7122,-0.379580), (7123,-0.542100), (7124,-0.585705), (7125,-0.742182), (7126,-0.486185), (7127,-0.642662), (7128,-0.960785), (7129,-1.115872), (7130,-0.471563), (7131,-0.619212), (7132,-0.651207), (7133,-0.838342), (7134,-0.869868), (7135,-0.989652), (7136,-1.040689), (7137,-1.221788), (7138,-0.555181), (7139,-0.713982), (7140,-0.787317), (7141,-0.913600), (7142,-0.695692), (7143,-0.835451), (7144,-0.903677), (7145,-1.046679), (7146,-0.376823), (7147,-0.539343), (7148,-0.601989), (7149,-0.715274), (7150,-0.748659), (7151,-0.867974), (7152,-0.915761), (7153,-1.040655), (7154,-0.395413), (7155,-0.531922), (7156,-0.600141), (7157,-0.745936), (7158,-0.505273), (7159,-0.682652), (7160,-0.644505), (7161,-0.810738), (7162,-0.510621), (7163,-0.247197), (7164,-0.308453), (7165,-0.449139), (7166,-0.427246), (7167,-0.603235), (7168,-0.750883), (7169,-0.885996), (7170,-0.627218), (7171,-0.387482), (7172,-0.413435), (7173,-0.593137), (7174,-0.456055), (7175,-0.501056), (7176,-0.729067), (7177,-0.884148), (7178,-0.609115), (7179,-0.367519), (7180,-0.391149), (7181,-0.541127), (7182,-0.483938), (7183,-0.695687), (7184,-0.717463), (7185,-0.895775), (7186,-0.622126), (7187,-0.394005), (7188,-0.473377), (7189,-0.615922), (7190,-0.448183), (7191,-0.519658), (7192,-0.761138), (7193,-0.491208), (7194,-0.631430), (7195,-0.277425), (7196,-0.454341), (7197,-0.458465), (7198,-0.601474), (7199,-0.684095), (7200,-0.818281), (7201,-0.537205), (7202,-0.647697), (7203,-0.340141), (7204,-0.500801), (7205,-0.351177), (7206,-0.515551), (7207,-0.471367), (7208,-0.927446), (7209,-0.636152), (7210,-0.412208), (7211,-0.448843), (7212,-0.592315), (7213,-0.601549), (7214,-0.775678), (7215,-0.824393), (7216,-0.971584), (7217,-0.678893), (7218,-0.486069), (7219,-0.533394), (7220,-0.698230), (7221,-0.532351), (7222,-0.594070), (7223,-0.639535), (7224,-0.747703), (7225,-0.471737), (7226,-0.607777), (7227,-0.282575), (7228,-0.445095), (7229,-0.430172), (7230,-0.603375), (7231,-0.664631), (7232,-0.831327), (7233,-0.533990), (7234,-0.678395), (7235,-0.351797), (7236,-0.518957), (7237,-0.399527), (7238,-0.532316), (7239,-0.505784), (7240,-0.730539), (7241,-0.471761), (7242,-0.605477), (7243,-0.312786), (7244,-0.463227), (7245,-0.456207), (7246,-0.584813), (7247,-0.656289), (7248,-0.825772), (7249,-0.571170), (7250,-0.695601), (7251,-0.374576), (7252,-0.520834), (7253,-0.444140), (7254,-0.603404), (7255,-0.547604), (7256,-0.776548), (7257,-0.520550), (7258,-0.682137), (7259,-0.309560), (7260,-0.484616), (7261,-0.481308), (7262,-0.573221), (7263,-0.680000), (7264,-0.829508), (7265,-0.551219), (7266,-0.691905), (7267,-0.368093), (7268,-0.536186), (7269,-0.356368), (7270,-0.517492), (7271,-0.497459), (7272,-0.876433), (7273,-0.607436), (7274,-0.315208), (7275,-0.377397), (7276,-0.514827), (7277,-0.514769), (7278,-0.689361), (7279,-0.739935), (7280,-0.914998), (7281,-0.634385), (7282,-0.357023), (7283,-0.402950), (7284,-0.575690), (7285,-0.414450), (7286,-0.488248), (7287,-0.540682), (7288,-0.916863), (7289,-0.629751), (7290,-0.380259), (7291,-0.457307), (7292,-0.612858), (7293,-0.600258), (7294,-0.766955), (7295,-0.799877), (7296,-1.258743), (7297,-0.953510), (7298,-0.737931), (7299,-0.812656), (7300,-0.981676), (7301,-0.840411), (7302,-0.901667), (7303,-0.973143), (7304,-1.019534), (7305,-1.160689), (7306,-0.482003), (7307,-0.625939), (7308,-0.682086), (7309,-0.796760), (7310,-0.791593), (7311,-0.931815), (7312,-1.021405), (7313,-1.173700), (7314,-0.486192), (7315,-0.648712), (7316,-0.677915), (7317,-0.815814), (7318,-0.597442), (7319,-0.762749), (7320,-1.027453), (7321,-1.172322), (7322,-0.504782), (7323,-0.681698), (7324,-0.742954), (7325,-0.910583), (7326,-0.891477), (7327,-1.056321), (7328,-1.108748), (7329,-1.261049), (7330,-0.561462), (7331,-0.753243), (7332,-0.820535), (7333,-0.951928), (7334,-0.705693), (7335,-0.852878), (7336,-1.014002), (7337,-1.177912), (7338,-0.475538), (7339,-0.637595), (7340,-0.661688), (7341,-0.807483), (7342,-0.848765), (7343,-0.989914), (7344,-1.052103), (7345,-1.201611), (7346,-0.523859), (7347,-0.688696), (7348,-0.742989), (7349,-0.889711), (7350,-0.677376), (7351,-0.836646), (7352,-1.164982), (7353,-1.293595), (7354,-0.596794), (7355,-0.709609), (7356,-0.776902), (7357,-0.913411), (7358,-0.923108), (7359,-1.101877), (7360,-1.145488), (7361,-1.298246), (7362,-0.622354), (7363,-0.780684), (7364,-0.840551), (7365,-0.998888), (7366,-0.764725), (7367,-0.878466), (7368,-0.944832), (7369,-1.076232), (7370,-0.411478), (7371,-0.552164), (7372,-0.603201), (7373,-0.757362), (7374,-0.793071), (7375,-0.922141), (7376,-0.975501), (7377,-1.162636), (7378,-0.461189), (7379,-0.640428), (7380,-0.674283), (7381,-0.815432), (7382,-0.583128), (7383,-0.771190), (7384,-1.064228), (7385,-1.248576), (7386,-0.599621), (7387,-0.704077), (7388,-0.808996), (7389,-0.937139), (7390,-0.962166), (7391,-1.136758), (7392,-1.213806), (7393,-1.334517), (7394,-0.640973), (7395,-0.751928), (7396,-0.827123), (7397,-0.969198), (7398,-0.733645), (7399,-0.926816), (7400,-0.956488), (7401,-1.109246), (7402,-0.441250), (7403,-0.577752), (7404,-0.643191), (7405,-0.785267), (7406,-0.824695), (7407,-0.974204), (7408,-1.070763), (7409,-1.198443), (7410,-0.508612), (7411,-0.658584), (7412,-0.698475), (7413,-0.868421), (7414,-0.634728), (7415,-0.773554), (7416,-0.746088), (7417,-0.882134), (7418,-0.598266), (7419,-0.345994), (7420,-0.441620), (7421,-0.632468), (7422,-0.594327), (7423,-0.759627), (7424,-0.766538), (7425,-0.913730), (7426,-0.663775), (7427,-0.428678), (7428,-0.448595), (7429,-0.635730), (7430,-0.474033), (7431,-0.611463), (7432,-0.814859), (7433,-0.947648), (7434,-0.644738), (7435,-0.394320), (7436,-0.498312), (7437,-0.634815), (7438,-0.598063), (7439,-0.808886), (7440,-0.852027), (7441,-1.030803), (7442,-0.765982), (7443,-0.522997), (7444,-0.550809), (7445,-0.678489), (7446,-0.513536), (7447,-0.598017), (7448,-0.871544), (7449,-0.606724), (7450,-0.769244), (7451,-0.444969), (7452,-0.554071), (7453,-0.542397), (7454,-0.686802), (7455,-0.746199), (7456,-0.912432), (7457,-0.644825), (7458,-0.816631), (7459,-0.485387), (7460,-0.627933), (7461,-0.481095), (7462,-0.651974), (7463,-0.621259), (7464,-1.003019), (7465,-0.745631), (7466,-0.464092), (7467,-0.510947), (7468,-0.710624), (7469,-0.711499), (7470,-0.874939), (7471,-0.932019), (7472,-1.107538), (7473,-0.816243), (7474,-0.618310), (7475,-0.702791), (7476,-0.853696), (7477,-0.687816), (7478,-0.742103), (7479,-0.789427), (7480,-0.918967), (7481,-0.647641), (7482,-0.801332), (7483,-0.471947), (7484,-0.615419), (7485,-0.620941), (7486,-0.713781), (7487,-0.800585), (7488,-0.946843), (7489,-0.652299), (7490,-0.855225), (7491,-0.497044), (7492,-0.634479), (7493,-0.471380), (7494,-0.619498), (7495,-0.605971), (7496,-0.857670), (7497,-0.611434), (7498,-0.737718), (7499,-0.366994), (7500,-0.556915), (7501,-0.499726), (7502,-0.670605), (7503,-0.770878), (7504,-0.919923), (7505,-0.613299), (7506,-0.771637), (7507,-0.416241), (7508,-0.589907), (7509,-0.465367), (7510,-0.600010), (7511,-0.546540), (7512,-0.831213), (7513,-0.573831), (7514,-0.699188), (7515,-0.386986), (7516,-0.562975), (7517,-0.556417), (7518,-0.704536), (7519,-0.777401), (7520,-0.915300), (7521,-0.636548), (7522,-0.781410), (7523,-0.438093), (7524,-0.644739), (7525,-0.505334), (7526,-0.636727), (7527,-0.598116), (7528,-0.992881), (7529,-0.708086), (7530,-0.432584), (7531,-0.446927), (7532,-0.616411), (7533,-0.605207), (7534,-0.788159), (7535,-0.849885), (7536,-1.008216), (7537,-0.707635), (7538,-0.464649), (7539,-0.537051), (7540,-0.693065), (7541,-0.542978), (7542,-0.626995), (7543,-0.693361), (7544,-1.135039), (7545,-0.819586), (7546,-0.568705), (7547,-0.601164), (7548,-0.764141), (7549,-0.739931), (7550,-0.899195), (7551,-0.997145), (7552,-1.092778), (7553,-0.828884), (7554,-0.952851), (7555,-0.625790), (7556,-0.757647), (7557,-0.600596), (7558,-0.735702), (7559,-0.706847), (7560,-0.875403), (7561,-1.023058), (7562,-0.772170), (7563,-0.537543), (7564,-0.593227), (7565,-0.766893), (7566,-0.753366), (7567,-0.949793), (7568,-1.005470), (7569,-1.157771), (7570,-0.827460), (7571,-0.623490), (7572,-0.665699), (7573,-0.823109), (7574,-0.672552), (7575,-0.766325), (7576,-0.917230), (7577,-1.089036), (7578,-0.800991), (7579,-0.588662), (7580,-0.629944), (7581,-0.787818), (7582,-0.755243), (7583,-0.916366), (7584,-0.994811), (7585,-1.152679), (7586,-0.848842), (7587,-0.613752), (7588,-0.694983), (7589,-0.869112), (7590,-0.693013), (7591,-0.756593), (7592,-1.109549), (7593,-1.228400), (7594,-0.571086), (7595,-0.728027), (7596,-0.789753), (7597,-0.938798), (7598,-0.922015), (7599,-1.078029), (7600,-1.160186), (7601,-1.300409), (7602,-0.591072), (7603,-0.754049), (7604,-0.808343), (7605,-0.951345), (7606,-0.693964), (7607,-0.864373), (7608,-0.961860), (7609,-1.085827), (7610,-0.821470), (7611,-0.570588), (7612,-0.591895), (7613,-0.743726), (7614,-0.765503), (7615,-0.952637), (7616,-1.017143), (7617,-1.185236), (7618,-0.891155), (7619,-0.643986), (7620,-0.712675), (7621,-0.890981), (7622,-0.734394), (7623,-0.759420), (7624,-0.866662), (7625,-1.023603), (7626,-0.734631), (7627,-0.504181), (7628,-0.530604), (7629,-0.695904), (7630,-0.700956), (7631,-0.863939), (7632,-0.928445), (7633,-1.089569), (7634,-0.794098), (7635,-0.568757), (7636,-0.627227), (7637,-0.777668), (7638,-0.669384), (7639,-0.721817), (7640,-0.947035), (7641,-1.075179), (7642,-0.778775), (7643,-0.535789), (7644,-0.605404), (7645,-0.756772), (7646,-0.748825), (7647,-0.906692), (7648,-0.966558), (7649,-1.127212), (7650,-0.810370), (7651,-0.573421), (7652,-0.604953), (7653,-0.799057), (7654,-0.634567), (7655,-0.732053), (7656,-0.778444), (7657,-0.890333), (7658,-0.656169), (7659,-0.399715), (7660,-0.435887), (7661,-0.600260), (7662,-0.575118), (7663,-0.760399), (7664,-0.797035), (7665,-0.963731), (7666,-0.689625), (7667,-0.447102), (7668,-0.528333), (7669,-0.691774), (7670,-0.540296), (7671,-0.629886), (7672,-0.808192), (7673,-0.973499), (7674,-0.695673), (7675,-0.435499), (7676,-0.490255), (7677,-0.662062), (7678,-0.647602), (7679,-0.831023), (7680,-0.911321), (7681,-1.051080), (7682,-0.790443), (7683,-0.542341), (7684,-0.567367), (7685,-0.754038), (7686,-0.587695), (7687,-0.658238), (7688,-0.885785), (7689,-1.019965), (7690,-0.738426), (7691,-0.484288), (7692,-0.593853), (7693,-0.741971), (7694,-0.721475), (7695,-0.886318), (7696,-0.920167), (7697,-1.121234), (7698,-0.875462), (7699,-0.612965), (7700,-0.646350), (7701,-0.787969), (7702,-0.636948), (7703,-0.727472), (7704,-0.961055), (7705,-0.693912), (7706,-0.844817), (7707,-0.479665), (7708,-0.632430), (7709,-0.652347), (7710,-0.782343), (7711,-0.873330), (7712,-1.001474), (7713,-0.760811), (7714,-0.919612), (7715,-0.577685), (7716,-0.748095), (7717,-0.563637), (7718,-0.704786), (7719,-0.661528), (7720,-0.862602), (7721,-0.598708), (7722,-0.764478), (7723,-0.442989), (7724,-0.592504), (7725,-0.599415), (7726,-0.754496), (7727,-0.837117), (7728,-0.950865), (7729,-0.656784), (7730,-0.803969), (7731,-0.459726), (7732,-0.618057), (7733,-0.461006), (7734,-0.607728), (7735,-0.578409), (7736,-0.949017), (7737,-0.657259), (7738,-0.809554), (7739,-0.496431), (7740,-0.638044), (7741,-0.629626), (7742,-0.795859), (7743,-0.856183), (7744,-1.000588), (7745,-0.770607), (7746,-0.930798), (7747,-0.552641), (7748,-0.714692), (7749,-0.567860), (7750,-0.717832), (7751,-0.681080), (7752,-0.940212), (7753,-0.677715), (7754,-0.794712), (7755,-0.449536), (7756,-0.604154), (7757,-0.586914), (7758,-0.755933), (7759,-0.826476), (7760,-1.004324), (7761,-0.709774), (7762,-0.914097), (7763,-0.577743), (7764,-0.721215), (7765,-0.537684), (7766,-0.771737), (7767,-0.704329), (7768,-0.943949), (7769,-0.646148), (7770,-0.797986), (7771,-0.457919), (7772,-0.621359), (7773,-0.625947), (7774,-0.750378), (7775,-0.838572), (7776,-1.004805), (7777,-0.722803), (7778,-0.877884), (7779,-0.544323), (7780,-0.690581), (7781,-0.522842), (7782,-0.657491), (7783,-0.647678), (7784,-1.033614), (7785,-0.725601), (7786,-0.493297), (7787,-0.533652), (7788,-0.712421), (7789,-0.696571), (7790,-0.867451), (7791,-0.928244), (7792,-1.078679), (7793,-0.752087), (7794,-0.522570), (7795,-0.591722), (7796,-0.752383), (7797,-0.612977), (7798,-0.688166), (7799,-0.716442), (7800,-0.917045), (7801,-0.637366), (7802,-0.760400), (7803,-0.472819), (7804,-0.598176), (7805,-0.627848), (7806,-0.776430), (7807,-0.807962), (7808,-1.102853), (7809,-1.327151), (7810,-0.659148), (7811,-0.828168), (7812,-0.864346), (7813,-1.024073), (7814,-0.756467), (7815,-0.894366), (7816,-0.987669), (7817,-1.125568), (7818,-0.458498), (7819,-0.603367), (7820,-0.633033), (7821,-0.782078), (7822,-0.790849), (7823,-0.939894), (7824,-0.998827), (7825,-1.156701), (7826,-0.472442), (7827,-0.627066), (7828,-0.692036), (7829,-0.847587), (7830,-0.607851), (7831,-0.746676), (7832,-0.979333), (7833,-1.041516), (7834,-0.822218), (7835,-0.539283), (7836,-0.718058), (7837,-0.774205), (7838,-0.917677), (7839,-0.928765), (7840,-1.071774), (7841,-1.125597), (7842,-0.850564), (7843,-0.601073), (7844,-0.710638), (7845,-0.753316), (7846,-0.784378), (7847,-0.683526), (7848,-0.920359), (7849,-0.996944), (7850,-0.791115), (7851,-0.477992), (7852,-0.669304), (7853,-0.744035), (7854,-0.902366), (7855,-0.885589), (7856,-1.040207), (7857,-1.084745), (7858,-0.856624), (7859,-0.584834), (7860,-0.758037), (7861,-0.786313), (7862,-0.865684), (7863,-0.685403), (7864,-1.084815), (7865,-1.153497), (7866,-0.904012), (7867,-0.602961), (7868,-0.767798), (7869,-0.798397), (7870,-0.970667), (7871,-1.000802), (7872,-1.174005), (7873,-1.209714), (7874,-0.949076), (7875,-0.677287), (7876,-0.835624), (7877,-0.892234), (7878,-0.929339), (7879,-0.767636), (7880,-0.863269), (7881,-0.932421), (7882,-0.704764), (7883,-0.412073), (7884,-0.568550), (7885,-0.633989), (7886,-0.790930), (7887,-0.747673), (7888,-0.934344), (7889,-0.981668), (7890,-0.757261), (7891,-0.524024), (7892,-0.737170), (7893,-0.812365), (7894,-0.854110), (7895,-0.695663), (7896,-1.080672), (7897,-1.133569), (7898,-0.899406), (7899,-0.649914), (7900,-0.801746), (7901,-0.822126), (7902,-1.029699), (7903,-1.020355), (7904,-1.164290), (7905,-1.194426), (7906,-0.939361), (7907,-0.676864), (7908,-0.846347), (7909,-0.887165), (7910,-0.942385), (7911,-0.822955), (7912,-0.992438), (7913,-1.028146), (7914,-0.803276), (7915,-0.477611), (7916,-0.649880), (7917,-0.696734), (7918,-0.835097), (7919,-0.789053), (7920,-0.954360), (7921,-1.026762), (7922,-0.774484), (7923,-0.482262), (7924,-0.647099), (7925,-0.727403), (7926,-0.794233), (7927,-0.634389), (7928,-0.683567), (7929,-0.736464), (7930,-0.892941), (7931,-0.233304), (7932,-0.388391), (7933,-0.452434), (7934,-0.588010), (7935,-0.577269), (7936,-0.756038), (7937,-0.803826), (7938,-0.955657), (7939,-0.282088), (7940,-0.449247), (7941,-0.494248), (7942,-0.660475), (7943,-0.415636), (7944,-0.744904), (7945,-0.801515), (7946,-0.952883), (7947,-0.311823), (7948,-0.438107), (7949,-0.491004), (7950,-0.647482), (7951,-0.654856), (7952,-0.788109), (7953,-0.828001), (7954,-1.010489), (7955,-0.345742), (7956,-0.486891), (7957,-0.542111), (7958,-0.718094), (7959,-0.484400), (7960,-0.753751), (7961,-0.922301), (7962,-0.648194), (7963,-0.410318), (7964,-0.433948), (7965,-0.631765), (7966,-0.589441), (7967,-0.748705), (7968,-0.810424), (7969,-0.943677), (7970,-0.703478), (7971,-0.473961), (7972,-0.536150), (7973,-0.693554), (7974,-0.537430), (7975,-0.570353), (7976,-0.885219), (7977,-1.080713), (7978,-0.398784), (7979,-0.601247), (7980,-0.610939), (7981,-0.786001), (7982,-0.772011), (7983,-0.929878), (7984,-0.975343), (7985,-1.136466), (7986,-0.455458), (7987,-0.622624), (7988,-0.681094), (7989,-0.858009), (7990,-0.602945), (7991,-0.764995), (7992,-0.805813), (7993,-0.944176), (7994,-0.647308), (7995,-0.377379), (7996,-0.426093), (7997,-0.574211), (7998,-0.557434), (7999,-0.723661), (8000,-0.796070), (8001,-0.951620), (8002,-0.677044), (8003,-0.419193), (8004,-0.448866), (8005,-0.619275), (8006,-0.463151), (8007,-0.536017), (8008,-0.697604), (8009,-0.863837), (8010,-0.586011), (8011,-0.343025), (8012,-0.414501), (8013,-0.565405), (8014,-0.544909), (8015,-0.712539), (8016,-0.773326), (8017,-0.904262), (8018,-0.617607), (8019,-0.372761), (8020,-0.453992), (8021,-0.625335), (8022,-0.474784), (8023,-0.548113), (8024,-0.705523), (8025,-0.858281), (8026,-0.562810), (8027,-0.337006), (8028,-0.370392), (8029,-0.544058), (8030,-0.504983), (8031,-0.701410), (8032,-0.790537), (8033,-0.931686), (8034,-0.655251), (8035,-0.411338), (8036,-0.456802), (8037,-0.596555), (8038,-0.490130), (8039,-0.585763), (8040,-0.871369), (8041,-1.061753), (8042,-0.356593), (8043,-0.517253), (8044,-0.571077), (8045,-0.709440), (8046,-0.675938), (8047,-0.840775), (8048,-0.905287), (8049,-1.038540), (8050,-0.356605), (8051,-0.496357), (8052,-0.564120), (8053,-0.718274), (8054,-0.485971), (8055,-0.648484), (8056,-0.954065), (8057,-1.111939), (8058,-0.449051), (8059,-0.612492), (8060,-0.691863), (8061,-0.813970), (8062,-0.849679), (8063,-0.985719), (8064,-0.877434), (8065,-0.626089), (8066,-0.355695), (8067,-0.503350), (8068,-0.545095), (8069,-0.623076), (8070,-0.438149), (8071,-0.615991), (8072,-0.752030), (8073,-0.406854), (8074,-0.574947), (8075,-0.299908), (8076,-0.463818), (8077,-0.568273), (8078,-0.710349), (8079,-0.695896), (8080,-0.848660), (8081,-0.504874), (8082,-0.659961), (8083,-0.410933), (8084,-0.568807), (8085,-0.515794), (8086,-0.668095), (8087,-0.503142), (8088,-0.661009), (8089,-0.712516), (8090,-0.440263), (8091,-0.159188), (8092,-0.308696), (8093,-0.323966), (8094,-0.522253), (8095,-0.529628), (8096,-0.692142), (8097,-0.742252), (8098,-0.502053), (8099,-0.209362), (8100,-0.393710), (8101,-0.408980), (8102,-0.494394), (8103,-0.352666), (8104,-0.652204), (8105,-0.330722), (8106,-0.457005), (8107,-0.228415), (8108,-0.350059), (8109,-0.436400), (8110,-0.592877), (8111,-0.564485), (8112,-0.751156), (8113,-0.395761), (8114,-0.567104), (8115,-0.273949), (8116,-0.410452), (8117,-0.410394), (8118,-0.567805), (8119,-0.416321), (8120,-0.829201), (8121,-0.499353), (8122,-0.645612), (8123,-0.369646), (8124,-0.521014), (8125,-0.586446), (8126,-0.730388), (8127,-0.716861), (8128,-0.840359), (8129,-0.498432), (8130,-0.670238), (8131,-0.424929), (8132,-0.597199), (8133,-0.534436), (8134,-0.685804), (8135,-0.554758), (8136,-0.746076), (8137,-0.400899), (8138,-0.555054), (8139,-0.301386), (8140,-0.468082), (8141,-0.513077), (8142,-0.680707), (8143,-0.654637), (8144,-0.843162), (8145,-0.491486), (8146,-0.635422), (8147,-0.372461), (8148,-0.541017), (8149,-0.527491), (8150,-0.665853), (8151,-0.519015), (8152,-0.668523), (8153,-0.682404), (8154,-0.422230), (8155,-0.153696), (8156,-0.309241), (8157,-0.371893), (8158,-0.555315), (8159,-0.552471), (8160,-0.656456), (8161,-0.719572), (8162,-0.482159), (8163,-0.195048), (8164,-0.345946), (8165,-0.382124), (8166,-0.469855), (8167,-0.314194), (8168,-0.501792), (8169,-0.555616), (8170,-0.335855), (8171,-0.049670), (8172,-0.208007), (8173,-0.271580), (8174,-0.417845), (8175,-0.414537), (8176,-0.585873), (8177,-0.651776), (8178,-0.379529), (8179,-0.117495), (8180,-0.257248), (8181,-0.326406), (8182,-0.393699), (8183,-0.245001), (8184,-0.430283), (8185,-0.516153), (8186,-0.292209), (8187,0.006518), (8188,-0.166221), (8189,-0.205643), (8190,-0.383028), (8191,-0.361136), (8192,-0.565459), (8193,-0.617886), (8194,-0.408807), (8195,-0.100794), (8196,-0.285605), (8197,-0.306912), (8198,-0.376534), (8199,-0.238519), (8200,-0.555251), (8201,-0.596996), (8202,-0.391167), (8203,-0.092910), (8204,-0.247991), (8205,-0.289272), (8206,-0.483376), (8207,-0.454057), (8208,-0.616571), (8209,-0.653213), (8210,-0.433915), (8211,-0.124036), (8212,-0.275873), (8213,-0.344562), (8214,-0.424397), (8215,-0.296137), (8216,-0.565951), (8217,-0.709423), (8218,-0.056755), (8219,-0.181649), (8220,-0.237326), (8221,-0.399382), (8222,-0.384922), (8223,-0.553015), (8224,-0.613808), (8225,-0.766566), (8226,-0.079521), (8227,-0.242505), (8228,-0.274964), (8229,-0.395675), (8230,-0.142933), (8231,-0.312416), (8232,-0.502337), (8233,-0.625835), (8234,0.036126), (8235,-0.131034), (8236,-0.216448), (8237,-0.374315), (8238,-0.374264), (8239,-0.514480), (8240,-0.587815), (8241,-0.736859), (8242,-0.051674), (8243,-0.218834), (8244,-0.244324), (8245,-0.412417), (8246,-0.166175), (8247,-0.324049), (8248,-0.512574), (8249,-0.675094), (8250,-0.024279), (8251,-0.174257), (8252,-0.209032), (8253,-0.378985), (8254,-0.372884), (8255,-0.520539), (8256,-0.568790), (8257,-0.711799), (8258,-0.075386), (8259,-0.245795), (8260,-0.288937), (8261,-0.428696), (8262,-0.196856), (8263,-0.342181), (8264,-0.487049), (8265,-0.637954), (8266,0.010074), (8267,-0.173347), (8268,-0.233207), (8269,-0.361351), (8270,-0.378481), (8271,-0.550287), (8272,-0.553015), (8273,-0.712286), (8274,-0.080049), (8275,-0.251392), (8276,-0.308002), (8277,-0.454261), (8278,-0.227530), (8279,-0.363106), (8280,-0.531662), (8281,-0.693713), (8282,0.010984), (8283,-0.148750), (8284,-0.204897), (8285,-0.368807), (8286,-0.363176), (8287,-0.501069), (8288,-0.553502), (8289,-0.703944), (8290,-0.002033), (8291,-0.132037), (8292,-0.216517), (8293,-0.403189), (8294,-0.162056), (8295,-0.335722), (8296,-0.579062), (8297,-0.363940), (8298,-0.073109), (8299,-0.250494), (8300,-0.287593), (8301,-0.444540), (8302,-0.445872), (8303,-0.594917), (8304,-0.635272), (8305,-0.395536), (8306,-0.139081), (8307,-0.313210), (8308,-0.363315), (8309,-0.447802), (8310,-0.254045), (8311,-0.410059), (8312,-0.690562), (8313,-0.473581), (8314,-0.234314), (8315,-0.383359), (8316,-0.401879), (8317,-0.555571), (8318,-0.543903), (8319,-0.706417), (8320,-0.612071), (8321,-0.773195), (8322,-0.250118), (8323,-0.393120), (8324,-0.468315), (8325,-0.633152), (8326,-0.286116), (8327,-0.438880), (8328,-0.724486), (8329,-0.478250), (8330,-0.447998), (8331,-0.623987), (8332,-0.681061), (8333,-0.863086), (8334,-0.562969), (8335,-0.718513), (8336,-0.768624), (8337,-0.500090), (8338,-0.388092), (8339,-0.520876), (8340,-0.557054), (8341,-0.659186), (8342,-0.371142), (8343,-0.511364), (8344,-0.519202), (8345,-0.680789), (8346,-0.309601), (8347,-0.457720), (8348,-0.512007), (8349,-0.656875), (8350,-0.394841), (8351,-0.565251), (8352,-0.623257), (8353,-0.759297), (8354,-0.234830), (8355,-0.400594), (8356,-0.449777), (8357,-0.601609), (8358,-0.267578), (8359,-0.421733), (8360,-0.709198), (8361,-0.362168), (8362,-0.488452), (8363,-0.479102), (8364,-0.626293), (8365,-0.724243), (8366,-0.884440), (8367,-0.651203), (8368,-0.778420), (8369,-0.413732), (8370,-0.565100), (8371,-0.409440), (8372,-0.558948), (8373,-0.535672), (8374,-0.727446), (8375,-0.435225), (8376,-0.608891), (8377,-0.652496), (8378,-0.433661), (8379,-0.380654), (8380,-0.556173), (8381,-0.583986), (8382,-0.771584), (8383,-0.505837), (8384,-0.653955), (8385,-0.703133), (8386,-0.454574), (8387,-0.310059), (8388,-0.505553), (8389,-0.551944), (8390,-0.619243), (8391,-0.341881), (8392,-0.638175), (8393,-0.316223), (8394,-0.448543), (8395,-0.434090), (8396,-0.566416), (8397,-0.696883), (8398,-0.838958), (8399,-0.563456), (8400,-0.719006), (8401,-0.403554), (8402,-0.534954), (8403,-0.402511), (8404,-0.505577), (8405,-0.469289), (8406,-0.632736), (8407,-0.370702), (8408,-0.522070), (8409,-0.596331), (8410,-0.343590), (8411,-0.342605), (8412,-0.510228), (8413,-0.558943), (8414,-0.726572), (8415,-0.416693), (8416,-0.598255), (8417,-0.628854), (8418,-0.420245), (8419,-0.284089), (8420,-0.442426), (8421,-0.476739), (8422,-0.549610), (8423,-0.274571), (8424,-0.442194), (8425,-0.472793), (8426,-0.273007), (8427,-0.250657), (8428,-0.384837), (8429,-0.448416), (8430,-0.640661), (8431,-0.350293), (8432,-0.523032), (8433,-0.582892), (8434,-0.337119), (8435,-0.178203), (8436,-0.337003), (8437,-0.375498), (8438,-0.432108), (8439,-0.156612), (8440,-0.364648), (8441,-0.432404), (8442,-0.190815), (8443,-0.178678), (8444,-0.335155), (8445,-0.407557), (8446,-0.585869), (8447,-0.322909), (8448,-0.452449), (8449,-0.510449), (8450,-0.258640), (8451,-0.121088), (8452,-0.261774), (8453,-0.332323), (8454,-0.386610), (8455,-0.128295), (8456,-0.432486), (8457,-0.493742), (8458,-0.252609), (8459,-0.250698), (8460,-0.375585), (8461,-0.456353), (8462,-0.600752), (8463,-0.337791), (8464,-0.487769), (8465,-0.543453), (8466,-0.268877), (8467,-0.129471), (8468,-0.304064), (8469,-0.345815), (8470,-0.428899), (8471,-0.136215), (8472,-0.503573), (8473,-0.664227), (8474,-0.275858), (8475,-0.425366), (8476,-0.466184), (8477,-0.601297), (8478,-0.357378), (8479,-0.516179), (8480,-0.569539), (8481,-0.734845), (8482,-0.192721), (8483,-0.316681), (8484,-0.392339), (8485,-0.544634), (8486,-0.152082), (8487,-0.314596), (8488,-0.389790), (8489,-0.589004), (8490,-0.154179), (8491,-0.291145), (8492,-0.365870), (8493,-0.528854), (8494,-0.297014), (8495,-0.429803), (8496,-0.478981), (8497,-0.628026), (8498,-0.099376), (8499,-0.238672), (8500,-0.299928), (8501,-0.465228), (8502,-0.098687), (8503,-0.241226), (8504,-0.427434), (8505,-0.596917), (8506,-0.208541), (8507,-0.384067), (8508,-0.414203), (8509,-0.527018), (8510,-0.308183), (8511,-0.449795), (8512,-0.493870), (8513,-0.630836), (8514,-0.060377), (8515,-0.224757), (8516,-0.291123), (8517,-0.435985), (8518,-0.081053), (8519,-0.239390), (8520,-0.377289), (8521,-0.536553), (8522,-0.146324), (8523,-0.289796), (8524,-0.357089), (8525,-0.503347), (8526,-0.230631), (8527,-0.378749), (8528,-0.420500), (8529,-0.588587), (8530,-0.016738), (8531,-0.189007), (8532,-0.241441), (8533,-0.382590), (8534,-0.032304), (8535,-0.180422), (8536,-0.431658), (8537,-0.602994), (8538,-0.198363), (8539,-0.356237), (8540,-0.395196), (8541,-0.529382), (8542,-0.294755), (8543,-0.454482), (8544,-0.529208), (8545,-0.681972), (8546,-0.120342), (8547,-0.282856), (8548,-0.352008), (8549,-0.476902), (8550,-0.103391), (8551,-0.271015), (8552,-0.539902), (8553,-0.283447), (8554,-0.268987), (8555,-0.418032), (8556,-0.463033), (8557,-0.620907), (8558,-0.353300), (8559,-0.514887), (8560,-0.558955), (8561,-0.335011), (8562,-0.180284), (8563,-0.361376), (8564,-0.462118), (8565,-0.542416), (8566,-0.272950), (8567,-0.412708), (8568,-0.527846), (8569,-0.655990), (8570,-0.252286), (8571,-0.376253), (8572,-0.450978), (8573,-0.602346), (8574,-0.344958), (8575,-0.477748), (8576,-0.645841), (8577,-0.659715), (8578,-0.441813), (8579,-0.293116), (8580,-0.425442), (8581,-0.478339), (8582,-0.526583), (8583,-0.226003), (8584,-0.502786), (8585,-0.556146), (8586,-0.363322), (8587,-0.313566), (8588,-0.436599), (8589,-0.498319), (8590,-0.687777), (8591,-0.385800), (8592,-0.560392), (8593,-0.603997), (8594,-0.389809), (8595,-0.246220), (8596,-0.431502), (8597,-0.457918), (8598,-0.520101), (8599,-0.220910), (8600,-0.484688), (8601,-0.532475), (8602,-0.292276), (8603,-0.287108), (8604,-0.429184), (8605,-0.470935), (8606,-0.624163), (8607,-0.391860), (8608,-0.545081), (8609,-0.629562), (8610,-0.371247), (8611,-0.197008), (8612,-0.379034), (8613,-0.418919), (8614,-0.491790), (8615,-0.226507), (8616,-0.677940), (8617,-0.345770), (8618,-0.496211), (8619,-0.470142), (8620,-0.641015), (8621,-0.705991), (8622,-0.856426), (8623,-0.579533), (8624,-0.746693), (8625,-0.389907), (8626,-0.559854), (8627,-0.447386), (8628,-0.590858), (8629,-0.551790), (8630,-0.713377), (8631,-0.468995), (8632,-0.636618), (8633,-0.697411), (8634,-0.470217), (8635,-0.419527), (8636,-0.583907), (8637,-0.641907), (8638,-0.837407), (8639,-0.571654), (8640,-0.700731), (8641,-0.769883), (8642,-0.523178), (8643,-0.355438), (8644,-0.506343), (8645,-0.581068), (8646,-0.620496), (8647,-0.324092), (8648,-0.535841), (8649,-0.587811), (8650,-0.352722), (8651,-0.364273), (8652,-0.482667), (8653,-0.556928), (8654,-0.719442), (8655,-0.423965), (8656,-0.605063), (8657,-0.660283), (8658,-0.408468), (8659,-0.237016), (8660,-0.433900), (8661,-0.475188), (8662,-0.541554), (8663,-0.281379), (8664,-0.604612), (8665,-0.628242), (8666,-0.429845), (8667,-0.419105), (8668,-0.545388), (8669,-0.603858), (8670,-0.793316), (8671,-0.495058), (8672,-0.615306), (8673,-0.680739), (8674,-0.433107), (8675,-0.265367), (8676,-0.439960), (8677,-0.488211), (8678,-0.562472), (8679,-0.301371), (8680,-0.346836), (8681,-0.514459), (8682,-0.168356), (8683,-0.329016), (8684,-0.335928), (8685,-0.495655), (8686,-0.575026), (8687,-0.694347), (8688,-0.399333), (8689,-0.528873), (8690,-0.191592), (8691,-0.377331), (8692,-0.206342), (8693,-0.354460), (8694,-0.334427), (8695,-0.482545), (8696,-0.473664), (8697,-0.521915), (8698,-0.308654), (8699,-0.277475), (8700,-0.434879), (8701,-0.466875), (8702,-0.666552), (8703,-0.381756), (8704,-0.513156), (8705,-0.591131), (8706,-0.391344), (8707,-0.192948), (8708,-0.321555), (8709,-0.365159), (8710,-0.438494), (8711,-0.160669), (8712,-0.351053), (8713,-0.498708), (8714,-0.148885), (8715,-0.332770), (8716,-0.322957), (8717,-0.485477), (8718,-0.549519), (8719,-0.675803), (8720,-0.423995), (8721,-0.569783), (8722,-0.238082), (8723,-0.367152), (8724,-0.248185), (8725,-0.392121), (8726,-0.370234), (8727,-0.545754), (8728,-0.509935), (8729,-0.666876), (8730,-0.255276), (8731,-0.385743), (8732,-0.448395), (8733,-0.586294), (8734,-0.358167), (8735,-0.516505), (8736,-0.554536), (8737,-0.726343), (8738,-0.166566), (8739,-0.315148), (8740,-0.401952), (8741,-0.530095), (8742,-0.182132), (8743,-0.334433), (8744,-0.407299), (8745,-0.440691), (8746,-0.233002), (8747,-0.190677), (8748,-0.342509), (8749,-0.394942), (8750,-0.557919), (8751,-0.306574), (8752,-0.459332), (8753,-0.524771), (8754,-0.254842), (8755,-0.118692), (8756,-0.242653), (8757,-0.312269), (8758,-0.380494), (8759,-0.144471), (8760,-0.549456), (8761,-0.705933), (8762,-0.283187), (8763,-0.432696), (8764,-0.493952), (8765,-0.659259), (8766,-0.400474), (8767,-0.560671), (8768,-0.632147), (8769,-0.769113), (8770,-0.232104), (8771,-0.384399), (8772,-0.437296), (8773,-0.604919), (8774,-0.229555), (8775,-0.409257), (8776,-0.545760), (8777,-0.576822), (8778,-0.322691), (8779,-0.303121), (8780,-0.441954), (8781,-0.488345), (8782,-0.683839), (8783,-0.405549), (8784,-0.535089), (8785,-0.609814), (8786,-0.358933), (8787,-0.237179), (8788,-0.361603), (8789,-0.397312), (8790,-0.468324), (8791,-0.175633), (8792,-0.437087), (8793,-0.604253), (8794,-0.186611), (8795,-0.343558), (8796,-0.408064), (8797,-0.569188), (8798,-0.302044), (8799,-0.463168), (8800,-0.514668), (8801,-0.685548), (8802,-0.151319), (8803,-0.263671), (8804,-0.348151), (8805,-0.469332), (8806,-0.101858), (8807,-0.284346), (8808,-0.533722), (8809,-0.199698), (8810,-0.336664), (8811,-0.325460), (8812,-0.494016), (8813,-0.562705), (8814,-0.685739), (8815,-0.397694), (8816,-0.564391), (8817,-0.254981), (8818,-0.389631), (8819,-0.250689), (8820,-0.406703), (8821,-0.372738), (8822,-0.514813), (8823,-0.269968), (8824,-0.422732), (8825,-0.481665), (8826,-0.268404), (8827,-0.247908), (8828,-0.385343), (8829,-0.448923), (8830,-0.609113), (8831,-0.331757), (8832,-0.621546), (8833,-0.699521), (8834,-0.445389), (8835,-0.296692), (8836,-0.472681), (8837,-0.539510), (8838,-0.616558), (8839,-0.324800), (8840,-0.607619), (8841,-0.660516), (8842,-0.362716), (8843,-0.371487), (8844,-0.544219), (8845,-0.613841), (8846,-0.799580), (8847,-0.527327), (8848,-0.678231), (8849,-0.724629), (8850,-0.453302), (8851,-0.295782), (8852,-0.454583), (8853,-0.504230), (8854,-0.563163), (8855,-0.304379), (8856,-0.646659), (8857,-0.731140), (8858,-0.491867), (8859,-0.467658), (8860,-0.648287), (8861,-0.705367), (8862,-0.879496), (8863,-0.615602), (8864,-0.758611), (8865,-0.830086), (8866,-0.579204), (8867,-0.403099), (8868,-0.575375), (8869,-0.627802), (8870,-0.716466), (8871,-0.437714), (8872,-0.542169), (8873,-0.670776), (8874,-0.319094), (8875,-0.490436), (8876,-0.473196), (8877,-0.631527), (8878,-0.688144), (8879,-0.862736), (8880,-0.593270), (8881,-0.736279), (8882,-0.381346), (8883,-0.517386), (8884,-0.361725), (8885,-0.509380), (8886,-0.458227), (8887,-0.623997), (8888,-0.615579), (8889,-0.674513), (8890,-0.448245), (8891,-0.430999), (8892,-0.589800), (8893,-0.649666), (8894,-0.809393), (8895,-0.528781), (8896,-0.680619), (8897,-0.737229), (8898,-0.490060), (8899,-0.326034), (8900,-0.531284), (8901,-0.555383), (8902,-0.644510), (8903,-0.369007), (8904,-0.467890), (8905,-0.618325), (8906,-0.265716), (8907,-0.405475), (8908,-0.404027), (8909,-0.557718), (8910,-0.640339), (8911,-0.805176), (8912,-0.539429), (8913,-0.681041), (8914,-0.325182), (8915,-0.469124), (8916,-0.325073), (8917,-0.488983), (8918,-0.476383), (8919,-0.596167), (8920,-0.673215), (8921,-0.720069), (8922,-0.497522), (8923,-0.486781), (8924,-0.663234), (8925,-0.686400), (8926,-0.882364), (8927,-0.604075), (8928,-0.758229), (8929,-0.834814), (8930,-0.557451), (8931,-0.389249), (8932,-0.561982), (8933,-0.636713), (8934,-0.699359), (8935,-0.412711), (8936,-0.452133), (8937,-0.597001), (8938,-0.266690), (8939,-0.427344), (8940,-0.429146), (8941,-0.606994), (8942,-0.654782), (8943,-0.804290), (8944,-0.534360), (8945,-0.701057), (8946,-0.337302), (8947,-0.495639), (8948,-0.337186), (8949,-0.508992), (8950,-0.510330), (8951,-0.680277), (8952,-0.550164), (8953,-0.599341), (8954,-0.366111), (8955,-0.335396), (8956,-0.535536), (8957,-0.581464), (8958,-0.728655), (8959,-0.471268), (8960,-0.572937), (8961,-0.636980), (8962,-0.390738), (8963,-0.245296), (8964,-0.410596), (8965,-0.447701), (8966,-0.525683), (8967,-0.252033), (8968,-0.472148), (8969,-0.624913), (8970,-0.266267), (8971,-0.429708), (8972,-0.412004), (8973,-0.559190), (8974,-0.625092), (8975,-0.795971), (8976,-0.526505), (8977,-0.701097), (8978,-0.318301), (8979,-0.482205), (8980,-0.320508), (8981,-0.453761), (8982,-0.438838), (8983,-0.583706), (8984,-0.408998), (8985,-0.480473), (8986,-0.629055), (8987,-0.232783), (8988,-0.379974), (8989,-0.447267), (8990,-0.577270), (8991,-0.331498), (8992,-0.480073), (8993,-0.533903), (8994,-0.708496), (8995,-0.184023), (8996,-0.344683), (8997,-0.388751), (8998,-0.509925), (8999,-0.159639), (9000,-0.570197), (9001,-0.620307), (9002,-0.382894), (9003,-0.357288), (9004,-0.522125), (9005,-0.559694), (9006,-0.770516), (9007,-0.478295), (9008,-0.657070), (9009,-0.674664), (9010,-0.444214), (9011,-0.273688), (9012,-0.453390), (9013,-0.493282), (9014,-0.548038), (9015,-0.257670), (9016,-0.522838), (9017,-0.574345), (9018,-0.366656), (9019,-0.338264), (9020,-0.497528), (9021,-0.565753), (9022,-0.720841), (9023,-0.451838), (9024,-0.580445), (9025,-0.612440), (9026,-0.407544), (9027,-0.272315), (9028,-0.429726), (9029,-0.482153), (9030,-0.536910), (9031,-0.265590), (9032,-0.519612), (9033,-0.584118), (9034,-0.359247), (9035,-0.362902), (9036,-0.521239), (9037,-0.588532), (9038,-0.722255), (9039,-0.432350), (9040,-0.610199), (9041,-0.670985), (9042,-0.423353), (9043,-0.275125), (9044,-0.453901), (9045,-0.503541), (9046,-0.559225), (9047,-0.250742), (9048,-0.421621), (9049,-0.527467), (9050,-0.663976), (9051,-0.270028), (9052,-0.437187), (9053,-0.494261), (9054,-0.630770), (9055,-0.401716), (9056,-0.546578), (9057,-0.591116), (9058,-0.730869), (9059,-0.164129), (9060,-0.322467), (9061,-0.360035), (9062,-0.471923), (9063,-0.103986), (9064,-0.488062), (9065,-0.563721), (9066,-0.319802), (9067,-0.313244), (9068,-0.469258), (9069,-0.503570), (9070,-0.681882), (9071,-0.389191), (9072,-0.554035), (9073,-0.610181), (9074,-0.337465), (9075,-0.182731), (9076,-0.371726), (9077,-0.399538), (9078,-0.453362), (9079,-0.168567), (9080,-0.505738), (9081,-0.603687), (9082,-0.339800), (9083,-0.354137), (9084,-0.508762), (9085,-0.577450), (9086,-0.736714), (9087,-0.463071), (9088,-0.816954), (9089,-0.857309), (9090,-0.616183), (9091,-0.468882), (9092,-0.610958), (9093,-0.689402), (9094,-0.758091), (9095,-0.460290), (9096,-0.729178), (9097,-0.790897), (9098,-0.573922), (9099,-0.558999), (9100,-0.673674), (9101,-0.720534), (9102,-0.911846), (9103,-0.588504), (9104,-0.765883), (9105,-0.834572), (9106,-0.560465), (9107,-0.435456), (9108,-0.564995), (9109,-0.628105), (9110,-0.709799), (9111,-0.450095), (9112,-0.431922), (9113,-0.613947), (9114,-0.675203), (9115,-0.442437), (9116,-0.409398), (9117,-0.559370), (9118,-0.606694), (9119,-0.806834), (9120,-0.525295), (9121,-0.722186), (9122,-0.772290), (9123,-0.506079), (9124,-0.348559), (9125,-0.519439), (9126,-0.566756), (9127,-0.631732), (9128,-0.534130), (9129,-0.663669), (9130,-0.323133), (9131,-0.459179), (9132,-0.469803), (9133,-0.622567), (9134,-0.689860), (9135,-0.847734), (9136,-0.581054), (9137,-0.715234), (9138,-0.363558), (9139,-0.515852), (9140,-0.362978), (9141,-0.582630), (9142,-0.544945), (9143,-0.669839), (9144,-0.690682), (9145,-0.843910), (9146,-0.517312), (9147,-0.672863), (9148,-0.658873), (9149,-0.833465), (9150,-0.863601), (9151,-1.017756), (9152,-0.729711), (9153,-0.866220), (9154,-0.534512), (9155,-0.677984), (9156,-0.528360), (9157,-0.673692), (9158,-0.629971), (9159,-0.787375), (9160,-0.553212), (9161,-0.711549), (9162,-0.377525), (9163,-0.548862), (9164,-0.516293), (9165,-0.675557), (9166,-0.729844), (9167,-0.849165), (9168,-0.606642), (9169,-0.764980), (9170,-0.402151), (9171,-0.540514), (9172,-0.405292), (9173,-0.545971), (9174,-0.517115), (9175,-0.691714), (9176,-0.428284), (9177,-0.581048), (9178,-0.640445), (9179,-0.393746), (9180,-0.379286), (9181,-0.556202), (9182,-0.590984), (9183,-0.743748), (9184,-0.468709), (9185,-0.637728), (9186,-0.686442), (9187,-0.467608), (9188,-0.315660), (9189,-0.464705), (9190,-0.527821), (9191,-0.592797), (9192,-0.347482), (9193,-0.487241), (9194,-0.554070), (9195,-0.293432), (9196,-0.258077), (9197,-0.424304), (9198,-0.444684), (9199,-0.651330), (9200,-0.374438), (9201,-0.534165), (9202,-0.550362), (9203,-0.339430), (9204,-0.198628), (9205,-0.368111), (9206,-0.385241), (9207,-0.456717), (9208,-0.235096), (9209,-0.440345), (9210,-0.473731), (9211,-0.210770), (9212,-0.178202), (9213,-0.331430), (9214,-0.393613), (9215,-0.578888), (9216,-0.336365), (9217,-0.503062), (9218,-0.562465), (9219,-0.295321), (9220,-0.156842), (9221,-0.300784), (9222,-0.357394), (9223,-0.425150), (9224,-0.309902), (9225,-0.472416), (9226,-0.512771), (9227,-0.236805), (9228,-0.237680), (9229,-0.408553), (9230,-0.495357), (9231,-0.639762), (9232,-0.367046), (9233,-0.501225), (9234,-0.573164), (9235,-0.337148), (9236,-0.167548), (9237,-0.316130), (9238,-0.366704), (9239,-0.431673), (9240,-0.459023), (9241,-0.538394), (9242,-0.687439), (9243,-0.293960), (9244,-0.485271), (9245,-0.508907), (9246,-0.664922), (9247,-0.387096), (9248,-0.520812), (9249,-0.609476), (9250,-0.770593), (9251,-0.234511), (9252,-0.398421), (9253,-0.469896), (9254,-0.590144), (9255,-0.256120), (9256,-0.437675), (9257,-0.537954), (9258,-0.669811), (9259,-0.260997), (9260,-0.412835), (9261,-0.491273), (9262,-0.608734), (9263,-0.351346), (9264,-0.503647), (9265,-0.552825), (9266,-0.694437), (9267,-0.162074), (9268,-0.330624), (9269,-0.367266), (9270,-0.509342), (9271,-0.161379), (9272,-0.409828), (9273,-0.491059), (9274,-0.621525), (9275,-0.228967), (9276,-0.380805), (9277,-0.458316), (9278,-0.606434), (9279,-0.355546), (9280,-0.488799), (9281,-0.578859), (9282,-0.710716), (9283,-0.174634), (9284,-0.314856), (9285,-0.366820), (9286,-0.527480), (9287,-0.157220), (9288,-0.390803), (9289,-0.458096), (9290,-0.632695), (9291,-0.211802), (9292,-0.370603), (9293,-0.429536), (9294,-0.578581), (9295,-0.338845), (9296,-0.455379), (9297,-0.511526), (9298,-0.701447), (9299,-0.157932), (9300,-0.259601), (9301,-0.319925), (9302,-0.501487), (9303,-0.126586), (9304,-0.462824), (9305,-0.522684), (9306,-0.670802), (9307,-0.280103), (9308,-0.420789), (9309,-0.495514), (9310,-0.641772), (9311,-0.361630), (9312,-0.525540), (9313,-0.622093), (9314,-0.776717), (9315,-0.244811), (9316,-0.360882), (9317,-0.422139), (9318,-0.563288), (9319,-0.185131), (9320,-0.501857), (9321,-0.525494), (9322,-0.295044), (9323,-0.284766), (9324,-0.477011), (9325,-0.521548), (9326,-0.675703), (9327,-0.389054), (9328,-0.545995), (9329,-0.596106), (9330,-0.341968), (9331,-0.210458), (9332,-0.352540), (9333,-0.380816), (9334,-0.435103), (9335,-0.180508), (9336,-0.587810), (9337,-0.657425), (9338,-0.441384), (9339,-0.391157), (9340,-0.515587), (9341,-0.571271), (9342,-0.792312), (9343,-0.510310), (9344,-0.665391), (9345,-0.710856), (9346,-0.857114), (9347,-0.334037), (9348,-0.452425), (9349,-0.505322), (9350,-0.669696), (9351,-0.334738), (9352,-0.702096), (9353,-0.765676), (9354,-0.565889), (9355,-0.564898), (9356,-0.710230), (9357,-0.782632), (9358,-0.937719), (9359,-0.645961), (9360,-0.825200), (9361,-0.868341), (9362,-0.637891), (9363,-0.455287), (9364,-0.628489), (9365,-0.686496), (9366,-0.765867), (9367,-0.483858), (9368,-0.453150), (9369,-0.612877), (9370,-0.663914), (9371,-0.414422), (9372,-0.413438), (9373,-0.559696), (9374,-0.641854), (9375,-0.806234), (9376,-0.503787), (9377,-0.691848), (9378,-0.730813), (9379,-0.474352), (9380,-0.302436), (9381,-0.470059), (9382,-0.535499), (9383,-0.594895), (9384,-0.583228), (9385,-0.749925), (9386,-0.412644), (9387,-0.557976), (9388,-0.563027), (9389,-0.700457), (9390,-0.777511), (9391,-0.933519), (9392,-0.666382), (9393,-0.832615), (9394,-0.511127), (9395,-0.651349), (9396,-0.479427), (9397,-0.621503), (9398,-0.645139), (9399,-0.791861), (9400,-0.530760), (9401,-0.674232), (9402,-0.725732), (9403,-0.472991), (9404,-0.491048), (9405,-0.640093), (9406,-0.732006), (9407,-0.914964), (9408,-0.681265), (9409,-0.804299), (9410,-0.832575), (9411,-0.600271), (9412,-0.448793), (9413,-0.607124), (9414,-0.633547), (9415,-0.697590), (9416,-0.564221), (9417,-0.752288), (9418,-0.422904), (9419,-0.570089), (9420,-0.574677), (9421,-0.710253), (9422,-0.798917), (9423,-0.947035), (9424,-0.683605), (9425,-0.849838), (9426,-0.468432), (9427,-0.622586), (9428,-0.471572), (9429,-0.642915), (9430,-0.611273), (9431,-0.762177), (9432,-0.553562), (9433,-0.692851), (9434,-0.745285), (9435,-0.473958), (9436,-0.460432), (9437,-0.615519), (9438,-0.654477), (9439,-0.840222), (9440,-0.556354), (9441,-0.719801), (9442,-0.768984), (9443,-0.545504), (9444,-0.406098), (9445,-0.568612), (9446,-0.629868), (9447,-0.711563), (9448,-0.409122), (9449,-0.527047), (9450,-0.613851), (9451,-0.348567), (9452,-0.369880), (9453,-0.514279), (9454,-0.553237), (9455,-0.761743), (9456,-0.452333), (9457,-0.619957), (9458,-0.666348), (9459,-0.423362), (9460,-0.270951), (9461,-0.433001), (9462,-0.507263), (9463,-0.545295), (9464,-0.316241), (9465,-0.478761), (9466,-0.520506), (9467,-0.264515), (9468,-0.272353), (9469,-0.400496), (9470,-0.471045), (9471,-0.627986), (9472,-0.350160), (9473,-0.524289), (9474,-0.582296), (9475,-0.356029), (9476,-0.189686), (9477,-0.345700), (9478,-0.420425), (9479,-0.505832), (9480,-0.367823), (9481,-0.520582), (9482,-0.601813), (9483,-0.373692), (9484,-0.364342), (9485,-0.518033), (9486,-0.569540), (9487,-0.706506), (9488,-0.401742), (9489,-0.575408), (9490,-0.626909), (9491,-0.389496), (9492,-0.235225), (9493,-0.383343), (9494,-0.433448), (9495,-0.520251), (9496,-0.553174), (9497,-0.628368), (9498,-0.762548), (9499,-0.373246), (9500,-0.513931), (9501,-0.556146), (9502,-0.707514), (9503,-0.473814), (9504,-0.622396), (9505,-0.710596), (9506,-0.845239), (9507,-0.275713), (9508,-0.434514), (9509,-0.474405), (9510,-0.653174), (9511,-0.317290), (9512,-0.522077), (9513,-0.591692), (9514,-0.747707), (9515,-0.337966), (9516,-0.478188), (9517,-0.567779), (9518,-0.675947), (9519,-0.432962), (9520,-0.588506), (9521,-0.658128), (9522,-0.809033), (9523,-0.259012), (9524,-0.423385), (9525,-0.437729), (9526,-0.585378), (9527,-0.217910), (9528,-0.486327), (9529,-0.523432), (9530,-0.682696), (9531,-0.292931), (9532,-0.443835), (9533,-0.485580), (9534,-0.625802), (9535,-0.373524), (9536,-0.510027), (9537,-0.569430), (9538,-0.719865), (9539,-0.158698), (9540,-0.281269), (9541,-0.344848), (9542,-0.513405), (9543,-0.162192), (9544,-0.428750), (9545,-0.451459), (9546,-0.628838), (9547,-0.210732), (9548,-0.396940), (9549,-0.413607), (9550,-0.569151), (9551,-0.302941), (9552,-0.462205), (9553,-0.536003), (9554,-0.743113), (9555,-0.180550), (9556,-0.324955), (9557,-0.397357), (9558,-0.555231), (9559,-0.170105), (9560,-0.485441), (9561,-0.558776), (9562,-0.715254), (9563,-0.299008), (9564,-0.436907), (9565,-0.515351), (9566,-0.653250), (9567,-0.400503), (9568,-0.593217), (9569,-0.642394), (9570,-0.781683), (9571,-0.250247), (9572,-0.406261), (9573,-0.465658), (9574,-0.620745), (9575,-0.267673), (9576,-0.668005), (9577,-0.715329), (9578,-0.463051), (9579,-0.476468), (9580,-0.606465), (9581,-0.667721), (9582,-0.839527), (9583,-0.508290), (9584,-0.660121), (9585,-0.712555), (9586,-0.465386), (9587,-0.338523), (9588,-0.480598), (9589,-0.500978), (9590,-0.571527), (9591,-0.326681), (9592,-0.509170), (9593,-0.551385), (9594,-0.703216), (9595,-0.325059), (9596,-0.481537), (9597,-0.536294), (9598,-0.700667), (9599,-0.418195), (9600,-0.744677), (9601,-0.788288), (9602,-0.559234), (9603,-0.384062), (9604,-0.533571), (9605,-0.597613), (9606,-0.672808), (9607,-0.401952), (9608,-0.564002), (9609,-0.692145), (9610,-0.365084), (9611,-0.517848), (9612,-0.521967), (9613,-0.695169), (9614,-0.770358), (9615,-0.907330), (9616,-0.642510), (9617,-0.783659), (9618,-0.434769), (9619,-0.607502), (9620,-0.472743), (9621,-0.642690), (9622,-0.636595), (9623,-0.789360), (9624,-0.453939), (9625,-0.599734), (9626,-0.625224), (9627,-0.407316), (9628,-0.404935), (9629,-0.621337), (9630,-0.625925), (9631,-0.803304), (9632,-0.568677), (9633,-0.714472), (9634,-0.724633), (9635,-0.494190), (9636,-0.327840), (9637,-0.512189), (9638,-0.566945), (9639,-0.644920), (9640,-0.537099), (9641,-0.705655), (9642,-0.353516), (9643,-0.500238), (9644,-0.474169), (9645,-0.607422), (9646,-0.675177), (9647,-0.830728), (9648,-0.561268), (9649,-0.707527), (9650,-0.377679), (9651,-0.544839), (9652,-0.419366), (9653,-0.556338), (9654,-0.543275), (9655,-0.703935), (9656,-0.668574), (9657,-0.832020), (9658,-0.520751), (9659,-0.649821), (9660,-0.631185), (9661,-0.760261), (9662,-0.844279), (9663,-0.984964), (9664,-0.707138), (9665,-0.878012), (9666,-0.537481), (9667,-0.686526), (9668,-0.525293), (9669,-0.698495), (9670,-0.664061), (9671,-0.816362), (9672,-0.587771), (9673,-0.736353), (9674,-0.400006), (9675,-0.545331), (9676,-0.537377), (9677,-0.698501), (9678,-0.777409), (9679,-0.908339), (9680,-0.633306), (9681,-0.794423), (9682,-0.429278), (9683,-0.605724), (9684,-0.454246), (9685,-0.608864), (9686,-0.570723), (9687,-0.748102), (9688,-0.497214), (9689,-0.643472), (9690,-0.681973), (9691,-0.412044), (9692,-0.435210), (9693,-0.571250), (9694,-0.611141), (9695,-0.866090), (9696,-0.587800), (9697,-0.753570), (9698,-0.817150), (9699,-0.561622), (9700,-0.405491), (9701,-0.553146), (9702,-0.614403), (9703,-0.672872), (9704,-0.415485), (9705,-0.575212), (9706,-0.622073), (9707,-0.388373), (9708,-0.341402), (9709,-0.537829), (9710,-0.580038), (9711,-0.752777), (9712,-0.438258), (9713,-0.615637), (9714,-0.668997), (9715,-0.455735), (9716,-0.264308), (9717,-0.422182), (9718,-0.470896), (9719,-0.526110), (9720,-0.322140), (9721,-0.453540), (9722,-0.513400), (9723,-0.279700), (9724,-0.259210), (9725,-0.408718), (9726,-0.451860), (9727,-0.634812), (9728,-0.314720), (9729,-0.495355), (9730,-0.558464), (9731,-0.312229), (9732,-0.163068), (9733,-0.325581), (9734,-0.352931), (9735,-0.431839), (9736,-0.303586), (9737,-0.461916), (9738,-0.511564), (9739,-0.253713), (9740,-0.226247), (9741,-0.409669), (9742,-0.437945), (9743,-0.614397), (9744,-0.320779), (9745,-0.505128), (9746,-0.553842), (9747,-0.315965), (9748,-0.170054), (9749,-0.331178), (9750,-0.383612), (9751,-0.449977), (9752,-0.494045), (9753,-0.571557), (9754,-0.699700), (9755,-0.290430), (9756,-0.462236), (9757,-0.510950), (9758,-0.685542), (9759,-0.460202), (9760,-0.570700), (9761,-0.612445), (9762,-0.797256), (9763,-0.252815), (9764,-0.413006), (9765,-0.471939), (9766,-0.615874), (9767,-0.238651), (9768,-0.420212), (9769,-0.452671), (9770,-0.603106), (9771,-0.181293), (9772,-0.347520), (9773,-0.380442), (9774,-0.529494), (9775,-0.301830), (9776,-0.455521), (9777,-0.489840), (9778,-0.615660), (9779,-0.064249), (9780,-0.235122), (9781,-0.307994), (9782,-0.481660), (9783,-0.102577), (9784,-0.365885), (9785,-0.426214), (9786,-0.586874), (9787,-0.196639), (9788,-0.349867), (9789,-0.409727), (9790,-0.542053), (9791,-0.306030), (9792,-0.431857), (9793,-0.502862), (9794,-0.654230), (9795,-0.113502), (9796,-0.249548), (9797,-0.328449), (9798,-0.508158), (9799,-0.178310), (9800,-0.382627), (9801,-0.449926), (9802,-0.605007), (9803,-0.184121), (9804,-0.351744), (9805,-0.414396), (9806,-0.558795), (9807,-0.322309), (9808,-0.470427), (9809,-0.539116), (9810,-0.679338), (9811,-0.149292), (9812,-0.296477), (9813,-0.338692), (9814,-0.497956), (9815,-0.135591), (9816,-0.503419), (9817,-0.565602), (9818,-0.728586), (9819,-0.312339), (9820,-0.442806), (9821,-0.496166), (9822,-0.660076), (9823,-0.386897), (9824,-0.531295), (9825,-0.616239), (9826,-0.755998), (9827,-0.244067), (9828,-0.387539), (9829,-0.451119), (9830,-0.606206), (9831,-0.226190), (9832,-0.358516), (9833,-0.533109), (9834,-0.215340), (9835,-0.349520), (9836,-0.345279), (9837,-0.480391), (9838,-0.552800), (9839,-0.699522), (9840,-0.446317), (9841,-0.618123), (9842,-0.256221), (9843,-0.419668), (9844,-0.247283), (9845,-0.458105), (9846,-0.417177), (9847,-0.575978), (9848,-0.659062), (9849,-0.704527), (9850,-0.432274), (9851,-0.409924), (9852,-0.589626), (9853,-0.642987), (9854,-0.839407), (9855,-0.543003), (9856,-0.594973), (9857,-0.785358), (9858,-0.834535), (9859,-0.597122), (9860,-0.473515), (9861,-0.621627), (9862,-0.654086), (9863,-0.717202), (9864,-0.677201), (9865,-0.804875), (9866,-0.470851), (9867,-0.631041), (9868,-0.622161), (9869,-0.790717), (9870,-0.825499), (9871,-0.969898), (9872,-0.707864), (9873,-0.837867), (9874,-0.510342), (9875,-0.667283), (9876,-0.526951), (9877,-0.692251), (9878,-0.663859), (9879,-0.802691), (9880,-0.507677), (9881,-0.653472), (9882,-0.696150), (9883,-0.430403), (9884,-0.429882), (9885,-0.614693), (9886,-0.672230), (9887,-0.828708), (9888,-0.545315), (9889,-0.712012), (9890,-0.745398), (9891,-0.510771), (9892,-0.404809), (9893,-0.564073), (9894,-0.641585), (9895,-0.697268), (9896,-0.999599), (9897,-0.763113), (9898,-0.495043), (9899,-0.561408), (9900,-0.678869), (9901,-0.697390), (9902,-0.876628), (9903,-0.911410), (9904,-1.072997), (9905,-0.784026), (9906,-0.553582), (9907,-0.598577), (9908,-0.743909), (9909,-0.597534), (9910,-0.641608), (9911,-0.708901), (9912,-0.610372), (9913,-0.783574), (9914,-0.839251), (9915,-0.612057), (9916,-0.601317), (9917,-0.747576), (9918,-0.786077), (9919,-0.971815), (9920,-0.708391), (9921,-0.846290), (9922,-0.893608), (9923,-0.640867), (9924,-0.484279), (9925,-0.628215), (9926,-0.678789), (9927,-0.731216), (9928,-0.944831), (9929,-0.647494), (9930,-0.431916), (9931,-0.482483), (9932,-0.617596), (9933,-0.599893), (9934,-0.795387), (9935,-0.840381), (9936,-1.014510), (9937,-0.726472), (9938,-0.472334), (9939,-0.518262), (9940,-0.686818), (9941,-0.539980), (9942,-0.618888), (9943,-0.679681), (9944,-0.560250), (9945,-0.709759), (9946,-0.742681), (9947,-0.471824), (9948,-0.478272), (9949,-0.663547), (9950,-0.741059), (9951,-0.914725), (9952,-0.622967), (9953,-0.778974), (9954,-0.834658), (9955,-0.549406), (9956,-0.408604), (9957,-0.586916), (9958,-0.604046), (9959,-0.709429), (9960,-0.740954), (9961,-0.458952), (9962,-0.636331), (9963,-0.299514), (9964,-0.453205), (9965,-0.430392), (9966,-0.567822), (9967,-0.667631), (9968,-0.815286), (9969,-0.521205), (9970,-0.672573), (9971,-0.389638), (9972,-0.517781), (9973,-0.369083), (9974,-0.542286), (9975,-0.490206), (9976,-0.386104), (9977,-0.537009), (9978,-0.579680), (9979,-0.376180), (9980,-0.351965), (9981,-0.520985), (9982,-0.548334), (9983,-0.740578), (9984,-0.399585), (9985,-0.567208), (9986,-0.595954), (9987,-0.372936), (9988,-0.230281), (9989,-0.398368), (9990,-0.414108), (9991,-0.506021), (9992,-0.709875), (9993,-0.448774), (9994,-0.602465), (9995,-0.248929), (9996,-0.421199), (9997,-0.416031), (9998,-0.559503), (9999,-0.644911), (10000,-0.750299), (10001,-0.475723), (10002,-0.662858), (10003,-0.365527), (10004,-0.531754), (10005,-0.392349), (10006,-0.531181), (10007,-0.492106), (10008,-0.537101), (10009,-0.707980), (10010,-0.727897), (10011,-0.496984), (10012,-0.490890), (10013,-0.635295), (10014,-0.684935), (10015,-0.817262), (10016,-0.527827), (10017,-0.668976), (10018,-0.727909), (10019,-0.493282), (10020,-0.328793), (10021,-0.508958), (10022,-0.566501), (10023,-0.604533), (10024,-0.365724), (10025,-0.532884), (10026,-0.580671), (10027,-0.372989), (10028,-0.349243), (10029,-0.508970), (10030,-0.571153), (10031,-0.762934), (10032,-0.495797), (10033,-0.643445), (10034,-0.730713), (10035,-0.495623), (10036,-0.328816), (10037,-0.465319), (10038,-0.531685), (10039,-0.631494), (10040,-0.441921), (10041,-0.609087), (10042,-0.582085), (10043,-0.338172), (10044,-0.347400), (10045,-0.518743), (10046,-0.574426), (10047,-0.746696), (10048,-0.486058), (10049,-0.650902), (10050,-0.693573), (10051,-0.452447), (10052,-0.300036), (10053,-0.448154), (10054,-0.481540), (10055,-0.561838), (10056,-0.363441), (10057,-0.546400), (10058,-0.597437), (10059,-0.373029), (10060,-0.371575), (10061,-0.542918), (10062,-0.624612), (10063,-0.818716), (10064,-0.537177), (10065,-0.719202), (10066,-0.783245), (10067,-0.504956), (10068,-0.342789), (10069,-0.493694), (10070,-0.539622), (10071,-0.588336), (10072,-0.463796), (10073,-0.646284), (10074,-0.680133), (10075,-0.438544), (10076,-0.391104), (10077,-0.586604), (10078,-0.622313), (10079,-0.811770), (10080,-0.546487), (10081,-0.688562), (10082,-0.767934), (10083,-0.507296), (10084,-0.344666), (10085,-0.489065), (10086,-0.517811), (10087,-0.614370), (10088,-0.537669), (10089,-0.681142), (10090,-0.343398), (10091,-0.489193), (10092,-0.480312), (10093,-0.650722), (10094,-0.734739), (10095,-0.879602), (10096,-0.621750), (10097,-0.776838), (10098,-0.416796), (10099,-0.565378), (10100,-0.412967), (10101,-0.575018), (10102,-0.556851), (10103,-0.723078), (10104,-0.496817), (10105,-0.634710), (10106,-0.657883), (10107,-0.413500), (10108,-0.423661), (10109,-0.532763), (10110,-0.583337), (10111,-0.762106), (10112,-0.589257), (10113,-0.759673), (10114,-0.789346), (10115,-0.569578), (10116,-0.442251), (10117,-0.597339), (10118,-0.630724), (10119,-0.705450), (10120,-0.530278), (10121,-0.678859), (10122,-0.747085), (10123,-0.519891), (10124,-0.497535), (10125,-0.690243), (10126,-0.768224), (10127,-0.968827), (10128,-0.659418), (10129,-0.822864), (10130,-0.824666), (10131,-0.603972), (10132,-0.457134), (10133,-0.644269), (10134,-0.695306), (10135,-0.758422), (10136,-0.577214), (10137,-0.725795), (10138,-0.770796), (10139,-0.518981), (10140,-0.476187), (10141,-0.652640), (10142,-0.691135), (10143,-0.856905), (10144,-0.569793), (10145,-0.740203), (10146,-0.806105), (10147,-0.562656), (10148,-0.418604), (10149,-0.593197), (10150,-0.611717), (10151,-0.647426), (10152,-0.637155), (10153,-0.800132), (10154,-0.484223), (10155,-0.631871), (10156,-0.583511), (10157,-0.741379), (10158,-0.837938), (10159,-0.967008), (10160,-0.699408), (10161,-0.859599), (10162,-0.502813), (10163,-0.676473), (10164,-0.533818), (10165,-0.693545), (10166,-0.649361), (10167,-0.784937), (10168,-0.537305), (10169,-0.705861), (10170,-0.772690), (10171,-0.524132), (10172,-0.514318), (10173,-0.681478), (10174,-0.723229), (10175,-0.915010), (10176,-0.644153), (10177,-0.811313), (10178,-0.838193), (10179,-0.596140), (10180,-0.454875), (10181,-0.620175), (10182,-0.678182), (10183,-0.708781), (10184,-0.449540), (10185,-0.618090), (10186,-0.681206), (10187,-0.413599), (10188,-0.434449), (10189,-0.600676), (10190,-0.657755), (10191,-0.848140), (10192,-0.598648), (10193,-0.748626), (10194,-0.794554), (10195,-0.568287), (10196,-0.446996), (10197,-0.570963), (10198,-0.622927), (10199,-0.683257), (10200,-0.590764), (10201,-0.754674), (10202,-0.794566), (10203,-0.522313), (10204,-0.523651), (10205,-0.679665), (10206,-0.705155), (10207,-0.869992), (10208,-0.572197), (10209,-0.729602), (10210,-0.816869), (10211,-0.549262), (10212,-0.389419), (10213,-0.603034), (10214,-0.623878), (10215,-0.702785), (10216,-0.718519), (10217,-0.446736), (10218,-0.576733), (10219,-0.230630), (10220,-0.409869), (10221,-0.409347), (10222,-0.569075), (10223,-0.629404), (10224,-0.787741), (10225,-0.525708), (10226,-0.675685), (10227,-0.343051), (10228,-0.501852), (10229,-0.368019), (10230,-0.503596), (10231,-0.464984), (10232,-0.449598), (10233,-0.605612), (10234,-0.664082), (10235,-0.415053), (10236,-0.409422), (10237,-0.563577), (10238,-0.603468), (10239,-0.781780), (10240,-1.091074), (10241,-0.812785), (10242,-0.982268), (10243,-0.685864), (10244,-0.828409), (10245,-0.693650), (10246,-0.835726), (10247,-0.792475), (10248,-1.003297), (10249,-1.130977), (10250,-0.862907), (10251,-0.614342), (10252,-0.663526), (10253,-0.836722), (10254,-0.846420), (10255,-0.994075), (10256,-1.025600), (10257,-1.172792), (10258,-0.884284), (10259,-0.617604), (10260,-0.673287), (10261,-0.841843), (10262,-0.681073), (10263,-0.767408), (10264,-0.915526), (10265,-0.639560), (10266,-0.818798), (10267,-0.867513), (10268,-0.576218), (10269,-0.576160), (10270,-0.742393), (10271,-0.818051), (10272,-0.978242), (10273,-0.684624), (10274,-0.866186), (10275,-0.938594), (10276,-0.692816), (10277,-0.537619), (10278,-0.709888), (10279,-0.781827), (10280,-0.990332), (10281,-0.719476), (10282,-0.914507), (10283,-0.539600), (10284,-0.710016), (10285,-0.686733), (10286,-0.836242), (10287,-0.898431), (10288,-1.025178), (10289,-0.765930), (10290,-0.898720), (10291,-0.552154), (10292,-0.736032), (10293,-0.569689), (10294,-0.730350), (10295,-0.733078), (10296,-1.079071), (10297,-0.795673), (10298,-0.944254), (10299,-0.626949), (10300,-0.774597), (10301,-0.773612), (10302,-0.898969), (10303,-0.923069), (10304,-1.087442), (10305,-0.840274), (10306,-0.971667), (10307,-0.608839), (10308,-0.768103), (10309,-0.703951), (10310,-0.831161), (10311,-0.786514), (10312,-1.056797), (10313,-0.785471), (10314,-0.943345), (10315,-0.608387), (10316,-0.750000), (10317,-0.748552), (10318,-0.890164), (10319,-0.977895), (10320,-1.136232), (10321,-0.839364), (10322,-0.991659), (10323,-0.644160), (10324,-0.758834), (10325,-0.625002), (10326,-0.780553), (10327,-0.761916), (10328,-0.881700), (10329,-0.603411), (10330,-0.788686), (10331,-0.798847), (10332,-0.555861), (10333,-0.539085), (10334,-0.705781), (10335,-0.783293), (10336,-0.959282), (10337,-0.653122), (10338,-0.802167), (10339,-0.859710), (10340,-0.632516), (10341,-0.455484), (10342,-0.629150), (10343,-0.698302), (10344,-1.116292), (10345,-0.835680), (10346,-0.609876), (10347,-0.653018), (10348,-0.799739), (10349,-0.800151), (10350,-0.996572), (10351,-1.017422), (10352,-1.176222), (10353,-0.882604), (10354,-0.635436), (10355,-0.712947), (10356,-0.879644), (10357,-0.720264), (10358,-0.797782), (10359,-0.840923), (10360,-1.018765), (10361,-0.711215), (10362,-0.894631), (10363,-0.548064), (10364,-0.708718), (10365,-0.688692), (10366,-0.832164), (10367,-0.934296), (10368,-1.292362), (10369,-0.996891), (10370,-0.771550), (10371,-0.797040), (10372,-0.966993), (10373,-0.817368), (10374,-0.897666), (10375,-0.960782), (10376,-1.207835), (10377,-0.953703), (10378,-0.691669), (10379,-0.787759), (10380,-0.940987), (10381,-0.936753), (10382,-1.144789), (10383,-1.184680), (10384,-1.317464), (10385,-1.078661), (10386,-0.825456), (10387,-0.867664), (10388,-1.035757), (10389,-0.866158), (10390,-0.895367), (10391,-0.951514), (10392,-1.178128), (10393,-1.328569), (10394,-0.653603), (10395,-0.821690), (10396,-0.875514), (10397,-1.029668), (10398,-1.041225), (10399,-1.217678), (10400,-1.279861), (10401,-1.460959), (10402,-0.750226), (10403,-0.887662), (10404,-0.950308), (10405,-1.078452), (10406,-0.863800), (10407,-1.013308), (10408,-1.078748), (10409,-1.215714), (10410,-0.540748), (10411,-0.716736), (10412,-0.806790), (10413,-0.957695), (10414,-0.957637), (10415,-1.074635), (10416,-1.131708), (10417,-1.300264), (10418,-0.639694), (10419,-0.789672), (10420,-0.854641), (10421,-0.995790), (10422,-0.762097), (10423,-0.929720), (10424,-1.155871), (10425,-1.283551), (10426,-0.617877), (10427,-0.805012), (10428,-0.843970), (10429,-1.023673), (10430,-1.025011), (10431,-1.193567), (10432,-1.261323), (10433,-1.384357), (10434,-0.704281), (10435,-0.846357), (10436,-0.886249), (10437,-1.052482), (10438,-0.819715), (10439,-0.976656), (10440,-1.076002), (10441,-1.231546), (10442,-0.560300), (10443,-0.709345), (10444,-0.743194), (10445,-0.923365), (10446,-0.960927), (10447,-1.103473), (10448,-1.149864), (10449,-1.318420), (10450,-0.652740), (10451,-0.809687), (10452,-0.903917), (10453,-1.058078), (10454,-0.833671), (10455,-0.962278), (10456,-1.271571), (10457,-1.438268), (10458,-0.770734), (10459,-0.917919), (10460,-0.968030), (10461,-1.083631), (10462,-1.066855), (10463,-1.219619), (10464,-1.296204), (10465,-1.447572), (10466,-0.770746), (10467,-0.910962), (10468,-0.976401), (10469,-1.143561), (10470,-0.909404), (10471,-1.044974), (10472,-1.098804), (10473,-1.259921), (10474,-0.605857), (10475,-0.764657), (10476,-0.811981), (10477,-0.966599), (10478,-0.971187), (10479,-1.150426), (10480,-1.199610), (10481,-1.365837), (10482,-0.691334), (10483,-0.856640), (10484,-0.910464), (10485,-1.034425), (10486,-0.764965), (10487,-0.912150), (10488,-0.849387), (10489,-1.019803), (10490,-0.770775), (10491,-0.530576), (10492,-0.589509), (10493,-0.701860), (10494,-0.719917), (10495,-0.920521), (10496,-0.926042), (10497,-1.068118), (10498,-0.794011), (10499,-0.562171), (10500,-0.623891), (10501,-0.786405), (10502,-0.643750), (10503,-0.707329), (10504,-0.927907), (10505,-1.073239), (10506,-0.810742), (10507,-0.567293), (10508,-0.621116), (10509,-0.766911), (10510,-0.785895), (10511,-0.966060), (10512,-1.024530), (10513,-1.173582), (10514,-0.906438), (10515,-0.698286), (10516,-0.730745), (10517,-0.887686), (10518,-0.701831), (10519,-0.780739), (10520,-1.035224), (10521,-0.761581), (10522,-0.906913), (10523,-0.573346), (10524,-0.701026), (10525,-0.702364), (10526,-0.843977), (10527,-0.910806), (10528,-1.084472), (10529,-0.785281), (10530,-0.941295), (10531,-0.598905), (10532,-0.746560), (10533,-0.609478), (10534,-0.750627), (10535,-0.745459), (10536,-1.137902), (10537,-0.848461), (10538,-0.625913), (10539,-0.687169), (10540,-0.839470), (10541,-0.851021), (10542,-1.021437), (10543,-1.067365), (10544,-1.219660), (10545,-0.936724), (10546,-0.723932), (10547,-0.765677), (10548,-0.899400), (10549,-0.722832), (10550,-0.824964), (10551,-0.870428), (10552,-1.023193), (10553,-0.743507), (10554,-0.893015), (10555,-0.560845), (10556,-0.697817), (10557,-0.673144), (10558,-0.834731), (10559,-0.914566), (10560,-1.102164), (10561,-0.795541), (10562,-0.947372), (10563,-0.602196), (10564,-0.769826), (10565,-0.621591), (10566,-0.764137), (10567,-0.734818), (10568,-0.979084), (10569,-0.709154), (10570,-0.838231), (10571,-0.529748), (10572,-0.687152), (10573,-0.667589), (10574,-0.825926), (10575,-0.894145), (10576,-1.055269), (10577,-0.815070), (10578,-0.950182), (10579,-0.577135), (10580,-0.737332), (10581,-0.590494), (10582,-0.713992), (10583,-0.680953), (10584,-0.938695), (10585,-0.654363), (10586,-0.827102), (10587,-0.480529), (10588,-0.630044), (10589,-0.601652), (10590,-0.770202), (10591,-0.842610), (10592,-1.009770), (10593,-0.744486), (10594,-0.930231), (10595,-0.586445), (10596,-0.726667), (10597,-0.590048), (10598,-0.719118), (10599,-0.706988), (10600,-1.084102), (10601,-0.810922), (10602,-0.586051), (10603,-0.638478), (10604,-0.780560), (10605,-0.778179), (10606,-0.952309), (10607,-1.001949), (10608,-1.131489), (10609,-0.857383), (10610,-0.621360), (10611,-0.691909), (10612,-0.855819), (10613,-0.713621), (10614,-0.770701), (10615,-0.822664), (10616,-1.123135), (10617,-0.833700), (10618,-0.629268), (10619,-0.676585), (10620,-0.861397), (10621,-0.838584), (10622,-1.014567), (10623,-1.047959), (10624,-1.295011), (10625,-1.029728), (10626,-0.780236), (10627,-0.865180), (10628,-1.016554), (10629,-0.858101), (10630,-0.917498), (10631,-0.970395), (10632,-1.240208), (10633,-0.944737), (10634,-0.701745), (10635,-0.789945), (10636,-0.943636), (10637,-0.925000), (10638,-1.094020), (10639,-1.131118), (10640,-1.289456), (10641,-1.013026), (10642,-0.757035), (10643,-0.818291), (10644,-0.981268), (10645,-0.829321), (10646,-0.916594), (10647,-0.992710), (10648,-1.341953), (10649,-1.056237), (10650,-0.813708), (10651,-0.844777), (10652,-0.998005), (10653,-0.964503), (10654,-1.165107), (10655,-1.209638), (10656,-1.351257), (10657,-1.082723), (10658,-0.879681), (10659,-0.918639), (10660,-1.088586), (10661,-0.903664), (10662,-0.964457), (10663,-1.024317), (10664,-1.086037), (10665,-1.255056), (10666,-0.602388), (10667,-0.732855), (10668,-0.803397), (10669,-0.964057), (10670,-0.966322), (10671,-1.130232), (10672,-1.184519), (10673,-1.339144), (10674,-0.639093), (10675,-0.780705), (10676,-0.834066), (10677,-0.978934), (10678,-0.733619), (10679,-0.885920), (10680,-1.247242), (10681,-0.959197), (10682,-0.728284), (10683,-0.764925), (10684,-0.929762), (10685,-0.919022), (10686,-1.088505), (10687,-1.170199), (10688,-1.346188), (10689,-1.053497), (10690,-0.831876), (10691,-0.881523), (10692,-1.027318), (10693,-0.874438), (10694,-0.964961), (10695,-1.020175), (10696,-1.121381), (10697,-1.227696), (10698,-0.527176), (10699,-0.677617), (10700,-0.767208), (10701,-0.930191), (10702,-0.932456), (10703,-1.063849), (10704,-1.122783), (10705,-1.306204), (10706,-0.644243), (10707,-0.793288), (10708,-0.881482), (10709,-1.016595), (10710,-0.792188), (10711,-0.956098), (10712,-1.329492), (10713,-1.014510), (10714,-0.787779), (10715,-0.842072), (10716,-1.014805), (10717,-1.018930), (10718,-1.209778), (10719,-1.239914), (10720,-1.414043), (10721,-1.110669), (10722,-0.864897), (10723,-0.927550), (10724,-1.090527), (10725,-0.924184), (10726,-1.000299), (10727,-1.078744), (10728,-1.132104), (10729,-1.278826), (10730,-0.569953), (10731,-0.730613), (10732,-0.779327), (10733,-0.926049), (10734,-0.957111), (10735,-1.101517), (10736,-1.144658), (10737,-1.322037), (10738,-0.686551), (10739,-0.808194), (10740,-0.847153), (10741,-0.999917), (10742,-0.762035), (10743,-0.916659), (10744,-0.978378), (10745,-0.711235), (10746,-0.857493), (10747,-0.532292), (10748,-0.664618), (10749,-0.661310), (10750,-0.811282), (10751,-0.903659), (10752,-1.079184), (10753,-0.806468), (10754,-0.929502), (10755,-0.559711), (10756,-0.713396), (10757,-0.580496), (10758,-0.727218), (10759,-0.721587), (10760,-0.962604), (10761,-1.108399), (10762,-0.786447), (10763,-0.584337), (10764,-0.640484), (10765,-0.781170), (10766,-0.750454), (10767,-0.931083), (10768,-0.978871), (10769,-1.120489), (10770,-0.877960), (10771,-0.630798), (10772,-0.652568), (10773,-0.826234), (10774,-0.672427), (10775,-0.749482), (10776,-1.024868), (10777,-0.749365), (10778,-0.877509), (10779,-0.518400), (10780,-0.703212), (10781,-0.671100), (10782,-0.854985), (10783,-0.946899), (10784,-1.125211), (10785,-0.845525), (10786,-0.994570), (10787,-0.630815), (10788,-0.810517), (10789,-0.642315), (10790,-0.773245), (10791,-0.743463), (10792,-1.153550), (10793,-0.877121), (10794,-0.629489), (10795,-0.693068), (10796,-0.868124), (10797,-0.853670), (10798,-1.017117), (10799,-1.110421), (10800,-1.261325), (10801,-0.979323), (10802,-0.746550), (10803,-0.761357), (10804,-0.903903), (10805,-0.754742), (10806,-0.809962), (10807,-0.900015), (10808,-1.034665), (10809,-0.748943), (10810,-0.926785), (10811,-0.614126), (10812,-0.747842), (10813,-0.728742), (10814,-0.914481), (10815,-0.951122), (10816,-1.095521), (10817,-0.836274), (10818,-0.977892), (10819,-0.633643), (10820,-0.774328), (10821,-0.614485), (10822,-0.783504), (10823,-0.722602), (10824,-0.967331), (10825,-0.684396), (10826,-0.831118), (10827,-0.491521), (10828,-0.618268), (10829,-0.631215), (10830,-0.798845), (10831,-0.892148), (10832,-1.039803), (10833,-0.766160), (10834,-0.948649), (10835,-0.624837), (10836,-0.795717), (10837,-0.615898), (10838,-0.744975), (10839,-0.736558), (10840,-0.986397), (10841,-0.730869), (10842,-0.852506), (10843,-0.481319), (10844,-0.669380), (10845,-0.655853), (10846,-0.823946), (10847,-0.901928), (10848,-1.021242), (10849,-0.758281), (10850,-0.906400), (10851,-0.562150), (10852,-0.730706), (10853,-0.578759), (10854,-0.731523), (10855,-0.698948), (10856,-1.044942), (10857,-0.801493), (10858,-0.552464), (10859,-0.584923), (10860,-0.744650), (10861,-0.716728), (10862,-0.899680), (10863,-0.983234), (10864,-1.147144), (10865,-0.851666), (10866,-0.614717), (10867,-0.647176), (10868,-0.792508), (10869,-0.657742), (10870,-0.734797), (10871,-0.801626), (10872,-1.096524), (10873,-0.844709), (10874,-0.616119), (10875,-0.697350), (10876,-0.831999), (10877,-0.767840), (10878,-0.958688), (10879,-1.018554), (10880,-1.374297), (10881,-1.109946), (10882,-0.867424), (10883,-0.912888), (10884,-1.070756), (10885,-0.921595), (10886,-1.005612), (10887,-1.039468), (10888,-1.183866), (10889,-1.346850), (10890,-0.674670), (10891,-0.803277), (10892,-0.842699), (10893,-0.975025), (10894,-1.007484), (10895,-1.094751), (10896,-1.146252), (10897,-1.305979), (10898,-0.629160), (10899,-0.808862), (10900,-0.867795), (10901,-1.040528), (10902,-0.798932), (10903,-0.936368), (10904,-1.100278), (10905,-1.259542), (10906,-0.562741), (10907,-0.746163), (10908,-0.801846), (10909,-0.968079), (10910,-0.959192), (10911,-1.096628), (10912,-1.137910), (10913,-1.291601), (10914,-0.635683), (10915,-0.787514), (10916,-0.819973), (10917,-0.981097), (10918,-0.737641), (10919,-0.905264), (10920,-1.229893), (10921,-1.009199), (10922,-0.747171), (10923,-0.926873), (10924,-0.985343), (10925,-1.135315), (10926,-1.135726), (10927,-1.287094), (10928,-1.339058), (10929,-1.087243), (10930,-0.831715), (10931,-0.983083), (10932,-1.008110), (10933,-1.087951), (10934,-0.923461), (10935,-1.094804), (10936,-1.177425), (10937,-1.336689), (10938,-0.683087), (10939,-0.822846), (10940,-0.891535), (10941,-1.054976), (10942,-1.052601), (10943,-1.206755), (10944,-1.272194), (10945,-1.419843), (10946,-0.771351), (10947,-0.911573), (10948,-0.940313), (10949,-1.106546), (10950,-0.870529), (10951,-1.000063), (10952,-1.101732), (10953,-1.242881), (10954,-0.602285), (10955,-0.779664), (10956,-0.809800), (10957,-0.950486), (10958,-0.970402), (10959,-1.117594), (10960,-1.209038), (10961,-1.329755), (10962,-0.651533), (10963,-0.785719), (10964,-0.855798), (10965,-1.000196), (10966,-0.810165), (10967,-0.965247), (10968,-1.188611), (10969,-1.320474), (10970,-0.625997), (10971,-0.735562), (10972,-0.826542), (10973,-0.956545), (10974,-0.979712), (10975,-1.132476), (10976,-1.179800), (10977,-1.339528), (10978,-0.705438), (10979,-0.821966), (10980,-0.845602), (10981,-1.008116), (10982,-0.769770), (10983,-0.919284), (10984,-0.987973), (10985,-1.136092), (10986,-0.486667), (10987,-0.645931), (10988,-0.689542), (10989,-0.859488), (10990,-0.865003), (10991,-1.019157), (10992,-1.072987), (10993,-1.200661), (10994,-0.516872), (10995,-0.688678), (10996,-0.727173), (10997,-0.870182), (10998,-0.665749), (10999,-0.805039), (11000,-0.997283), (11001,-1.148651), (11002,-0.477398), (11003,-0.647814), (11004,-0.726252), (11005,-0.888309), (11006,-0.879422), (11007,-1.038223), (11008,-1.060926), (11009,-1.197898), (11010,-0.540114), (11011,-0.711920), (11012,-0.759708), (11013,-0.905503), (11014,-0.661120), (11015,-0.813422), (11016,-1.036323), (11017,-1.199300), (11018,-0.521084), (11019,-0.684061), (11020,-0.739745), (11021,-0.867425), (11022,-0.876196), (11023,-1.066580), (11024,-1.133873), (11025,-1.285241), (11026,-0.653474), (11027,-0.819244), (11028,-0.862848), (11029,-1.014216), (11030,-0.770297), (11031,-0.927238), (11032,-1.202631), (11033,-0.941994), (11034,-0.674850), (11035,-0.721705), (11036,-0.865640), (11037,-0.860479), (11038,-1.025316), (11039,-1.051269), (11040,-1.250946), (11041,-0.962437), (11042,-0.706909), (11043,-0.737972), (11044,-0.910711), (11045,-0.767586), (11046,-0.811197), (11047,-0.858052), (11048,-1.031248), (11049,-0.764111), (11050,-0.505327), (11051,-0.580985), (11052,-0.721670), (11053,-0.717899), (11054,-0.899924), (11055,-0.941669), (11056,-1.107439), (11057,-0.854698), (11058,-0.614961), (11059,-0.663212), (11060,-0.843378), (11061,-0.688180), (11062,-0.749900), (11063,-0.815339), (11064,-1.138108), (11065,-0.886293), (11066,-0.631692), (11067,-0.673443), (11068,-0.843853), (11069,-0.826143), (11070,-0.997023), (11071,-1.055029), (11072,-1.216616), (11073,-0.943436), (11074,-0.679079), (11075,-0.749628), (11076,-0.916788), (11077,-0.766700), (11078,-0.831206), (11079,-0.843227), (11080,-1.116297), (11081,-0.839398), (11082,-0.591303), (11083,-0.666954), (11084,-0.822969), (11085,-0.865183), (11086,-1.025374), (11087,-1.043437), (11088,-1.200378), (11089,-0.910943), (11090,-0.681889), (11091,-0.727354), (11092,-0.905659), (11093,-0.744426), (11094,-0.807072), (11095,-0.890627), (11096,-1.143722), (11097,-0.845921), (11098,-0.612691), (11099,-0.643753), (11100,-0.815096), (11101,-0.774162), (11102,-0.938072), (11103,-1.004438), (11104,-1.188323), (11105,-0.923502), (11106,-0.711174), (11107,-0.771967), (11108,-0.915902), (11109,-0.770454), (11110,-0.875373), (11111,-0.894363), (11112,-1.283550), (11113,-0.563994), (11114,-0.746019), (11115,-0.795660), (11116,-0.946565), (11117,-0.918179), (11118,-1.079296), (11119,-1.139626), (11120,-1.294244), (11121,-0.598839), (11122,-0.760427), (11123,-0.818896), (11124,-0.980947), (11125,-0.744467), (11126,-0.905121), (11127,-0.980316), (11128,-1.166054), (11129,-0.849675), (11130,-0.590897), (11131,-0.663769), (11132,-0.822100), (11133,-0.804860), (11134,-0.995708), (11135,-1.011448), (11136,-1.327247), (11137,-1.485115), (11138,-0.802716), (11139,-0.973132), (11140,-1.019060), (11141,-1.184360), (11142,-0.937661), (11143,-1.079737), (11144,-1.261299), (11145,-1.390369), (11146,-0.752096), (11147,-0.881636), (11148,-0.956825), (11149,-1.098907), (11150,-1.121146), (11151,-1.267868), (11152,-1.313796), (11153,-1.462841), (11154,-0.787411), (11155,-0.952248), (11156,-0.990743), (11157,-1.164409), (11158,-0.933032), (11159,-1.073718), (11160,-1.059728), (11161,-1.134916), (11162,-1.289540), (11163,-0.636402), (11164,-0.766869), (11165,-0.833235), (11166,-0.995285), (11167,-1.006843), (11168,-1.150778), (11169,-1.194383), (11170,-1.351323), (11171,-0.710734), (11172,-0.823549), (11173,-0.908956), (11174,-1.056148), (11175,-0.828948), (11176,-1.164722), (11177,-1.218082), (11178,-0.950475), (11179,-0.672656), (11180,-0.812409), (11181,-0.891780), (11182,-1.041758), (11183,-1.039377), (11184,-1.193994), (11185,-1.252464), (11186,-1.021094), (11187,-0.717720), (11188,-0.897422), (11189,-0.948923), (11190,-1.004143), (11191,-0.837794), (11192,-1.277149), (11193,-1.330046), (11194,-1.119577), (11195,-0.841288), (11196,-1.022843), (11197,-1.064594), (11198,-1.205743), (11199,-1.198716), (11200,-1.390497), (11201,-1.420633), (11202,-1.193439), (11203,-0.928155), (11204,-1.070700), (11205,-1.107336), (11206,-1.201572), (11207,-1.058454), (11208,-1.250228), (11209,-1.286870), (11210,-1.035518), (11211,-0.758162), (11212,-0.904421), (11213,-0.958244), (11214,-1.123081), (11215,-1.096086), (11216,-1.253026), (11217,-1.303600), (11218,-1.059681), (11219,-0.775356), (11220,-0.929047), (11221,-0.974511), (11222,-1.031585), (11223,-0.890326), (11224,-1.093253), (11225,-1.128498), (11226,-1.290549), (11227,-0.614186), (11228,-0.792961), (11229,-0.859791), (11230,-0.989794), (11231,-1.002741), (11232,-1.150396), (11233,-1.198184), (11234,-1.326790), (11235,-0.656001), (11236,-0.801796), (11237,-0.867235), (11238,-1.031145), (11239,-0.821597), (11240,-0.958569), (11241,-0.996601), (11242,-1.148895), (11243,-0.481362), (11244,-0.637839), (11245,-0.675871), (11246,-0.863006), (11247,-0.852729), (11248,-1.025931), (11249,-1.098797), (11250,-1.225550), (11251,-0.590527), (11252,-0.747005), (11253,-0.805011), (11254,-0.938264), (11255,-0.731045), (11256,-0.920503), (11257,-0.965967), (11258,-1.121512), (11259,-0.464661), (11260,-0.583981), (11261,-0.622013), (11262,-0.778491), (11263,-0.836960), (11264,-0.977176), (11265,-1.048188), (11266,-1.200020), (11267,-0.538992), (11268,-0.687104), (11269,-0.725605), (11270,-0.858395), (11271,-0.694369), (11272,-1.019461), (11273,-1.068638), (11274,-1.207927), (11275,-0.553863), (11276,-0.701518), (11277,-0.769743), (11278,-0.919715), (11279,-0.896432), (11280,-1.052446), (11281,-1.105807), (11282,-1.270180), (11283,-0.617512), (11284,-0.770733), (11285,-0.807375), (11286,-0.970358), (11287,-0.738982), (11288,-1.005076), (11289,-1.149945), (11290,-0.839608), (11291,-0.607298), (11292,-0.660195), (11293,-0.814819), (11294,-0.795713), (11295,-0.957300), (11296,-1.022276), (11297,-1.176894), (11298,-0.902324), (11299,-0.667698), (11300,-0.715479), (11301,-0.852915), (11302,-0.707473), (11303,-0.771053), (11304,-0.967937), (11305,-1.131847), (11306,-0.820584), (11307,-0.604535), (11308,-0.655109), (11309,-0.824129), (11310,-0.792017), (11311,-0.962897), (11312,-1.033909), (11313,-1.197356), (11314,-0.901415), (11315,-0.669111), (11316,-0.665804), (11317,-0.842719), (11318,-0.708887), (11319,-0.836567), (11320,-0.995367), (11321,-1.138370), (11322,-0.834539), (11323,-0.608272), (11324,-0.650950), (11325,-0.818573), (11326,-0.786931), (11327,-0.977316), (11328,-0.975868), (11329,-1.148601), (11330,-0.879140), (11331,-0.652410), (11332,-0.717379), (11333,-0.877576), (11334,-0.704264), (11335,-0.800354), (11336,-0.936393), (11337,-1.137930), (11338,-0.794144), (11339,-0.556267), (11340,-0.561782), (11341,-0.767032), (11342,-0.707989), (11343,-0.896514), (11344,-0.964739), (11345,-1.113321), (11346,-0.847574), (11347,-0.588790), (11348,-0.655156), (11349,-0.800487), (11350,-0.693136), (11351,-0.742313), (11352,-0.926198), (11353,-1.088248), (11354,-0.844329), (11355,-0.601344), (11356,-0.628693), (11357,-0.771702), (11358,-0.769784), (11359,-0.943450), (11360,-1.013065), (11361,-1.175116), (11362,-0.913088), (11363,-0.647804), (11364,-0.681653), (11365,-0.838131), (11366,-0.713128), (11367,-0.795285), (11368,-1.037228), (11369,-1.172804), (11370,-0.490406), (11371,-0.658035), (11372,-0.700244), (11373,-0.843716), (11374,-0.863169), (11375,-0.981557), (11376,-1.066501), (11377,-1.238307), (11378,-0.566127), (11379,-0.707746), (11380,-0.736022), (11381,-0.901322), (11382,-0.670878), (11383,-0.807845), (11384,-1.126431), (11385,-1.262007), (11386,-0.581931), (11387,-0.738872), (11388,-0.793629), (11389,-0.933851), (11390,-0.935183), (11391,-1.114891), (11392,-1.386559), (11393,-1.539323), (11394,-0.893154), (11395,-1.029194), (11396,-1.042611), (11397,-1.182827), (11398,-0.992326), (11399,-1.140444), (11400,-1.284380), (11401,-1.445040), (11402,-0.775184), (11403,-0.928875), (11404,-0.973406), (11405,-1.127567), (11406,-1.153520), (11407,-1.282127), (11408,-1.382863), (11409,-1.542133), (11410,-0.856015), (11411,-1.005060), (11412,-1.093260), (11413,-1.245555), (11414,-1.024397), (11415,-1.146968), (11416,-1.176177), (11417,-1.230464), (11418,-1.347461), (11419,-0.672025), (11420,-0.823863), (11421,-0.889766), (11422,-1.049030), (11423,-1.040612), (11424,-1.187797), (11425,-1.269955), (11426,-1.388813), (11427,-0.741711), (11428,-0.878220), (11429,-0.939940), (11430,-1.090375), (11431,-0.888728), (11432,-1.263519), (11433,-1.348000), (11434,-1.045559), (11435,-0.786782), (11436,-0.962764), (11437,-0.989187), (11438,-1.195363), (11439,-1.181373), (11440,-1.327632), (11441,-1.348012), (11442,-1.121281), (11443,-0.869003), (11444,-1.030127), (11445,-1.061659), (11446,-1.124305), (11447,-0.982577), (11448,-1.381988), (11449,-1.446495), (11450,-1.139408), (11451,-0.849973), (11452,-1.022242), (11453,-1.081639), (11454,-1.267384), (11455,-1.243631), (11456,-1.395469), (11457,-1.432568), (11458,-1.194691), (11459,-0.934981), (11460,-1.088672), (11461,-1.123917), (11462,-1.219550), (11463,-1.050414), (11464,-1.240799), (11465,-1.315530), (11466,-1.046990), (11467,-0.768701), (11468,-0.929825), (11469,-0.941382), (11470,-1.130377), (11471,-1.133105), (11472,-1.284936), (11473,-1.340157), (11474,-1.128755), (11475,-0.847679), (11476,-0.991151), (11477,-1.048224), (11478,-1.145711), (11479,-1.012348), (11480,-1.166966), (11481,-1.218936), (11482,-1.356366), (11483,-0.719489), (11484,-0.846236), (11485,-0.897273), (11486,-1.046788), (11487,-1.079247), (11488,-1.240364), (11489,-1.315559), (11490,-1.452525), (11491,-0.767803), (11492,-0.914995), (11493,-0.990647), (11494,-1.129479), (11495,-0.909248), (11496,-1.046684), (11497,-1.089825), (11498,-1.245376), (11499,-0.581556), (11500,-0.727351), (11501,-0.778851), (11502,-0.939505), (11503,-0.912973), (11504,-1.060628), (11505,-1.115848), (11506,-1.270002), (11507,-0.601536), (11508,-0.745471), (11509,-0.828562), (11510,-1.013373), (11511,-0.797789), (11512,-0.991893), (11513,-1.062441), (11514,-1.202194), (11515,-0.543483), (11516,-0.689741), (11517,-0.743571), (11518,-0.887044), (11519,-0.913460), (11520,-1.048109), (11521,-1.099146), (11522,-1.261660), (11523,-0.577865), (11524,-0.755250), (11525,-0.825793), (11526,-0.975307), (11527,-0.715596), (11528,-1.037432), (11529,-1.113554), (11530,-1.293256), (11531,-0.595528), (11532,-0.738537), (11533,-0.820695), (11534,-0.959521), (11535,-0.980834), (11536,-1.142884), (11537,-1.151655), (11538,-1.311383), (11539,-0.647562), (11540,-0.794284), (11541,-0.850894), (11542,-0.984153), (11543,-0.753240), (11544,-1.099697), (11545,-1.251528), (11546,-0.973702), (11547,-0.738612), (11548,-0.786400), (11549,-0.978644), (11550,-0.960934), (11551,-1.102083), (11552,-1.188887), (11553,-1.319354), (11554,-1.045711), (11555,-0.806901), (11556,-0.875590), (11557,-1.028355), (11558,-0.852256), (11559,-0.928841), (11560,-1.018431), (11561,-1.173512), (11562,-0.885468), (11563,-0.651774), (11564,-0.735328), (11565,-0.887160), (11566,-0.854585), (11567,-1.021751), (11568,-1.087184), (11569,-1.217187), (11570,-0.945404), (11571,-0.697765), (11572,-0.755308), (11573,-0.939193), (11574,-0.787246), (11575,-0.826668), (11576,-0.969676), (11577,-1.135446), (11578,-0.844615), (11579,-0.611385), (11580,-0.669385), (11581,-0.827722), (11582,-0.828134), (11583,-1.011086), (11584,-1.073732), (11585,-1.216277), (11586,-0.937525), (11587,-0.701039), (11588,-0.752076), (11589,-0.899731), (11590,-0.779367), (11591,-0.799284), (11592,-0.991528), (11593,-1.120605), (11594,-0.870186), (11595,-0.625804), (11596,-0.648507), (11597,-0.832855), (11598,-0.866241), (11599,-0.979519), (11600,-1.065396), (11601,-1.245562), (11602,-0.940798), (11603,-0.712208), (11604,-0.772537), (11605,-0.920656), (11606,-0.774281), (11607,-0.857366), (11608,-1.077017), (11609,-1.201447), (11610,-0.910616), (11611,-0.683422), (11612,-0.727954), (11613,-0.876998), (11614,-0.894129), (11615,-1.086373), (11616,-1.145306), (11617,-1.288778), (11618,-0.988198), (11619,-0.781435), (11620,-0.843625), (11621,-0.971768), (11622,-0.800309), (11623,-0.836488), (11624,-1.031518), (11625,-1.179637), (11626,-0.521389), (11627,-0.674147), (11628,-0.736336), (11629,-0.891418), (11630,-0.882537), (11631,-1.031118), (11632,-1.167158), (11633,-1.302734), (11634,-0.621732), (11635,-0.785172), (11636,-0.847825), (11637,-0.971785), (11638,-0.754810), (11639,-0.894106), (11640,-1.206186), (11641,-1.338976), (11642,-0.702563), (11643,-0.843248), (11644,-0.907754), (11645,-1.029862), (11646,-1.043736), (11647,-1.196037), (11648,-1.218740), (11649,-1.370108), (11650,-1.103898), (11651,-0.851619), (11652,-0.912876), (11653,-1.068890), (11654,-0.911833), (11655,-1.006996), (11656,-1.138853), (11657,-1.326457), (11658,-1.043058), (11659,-0.783811), (11660,-0.814873), (11661,-1.003868), (11662,-0.986158), (11663,-1.181189), (11664,-1.225263), (11665,-1.397069), (11666,-1.110421), (11667,-0.881367), (11668,-0.927758), (11669,-1.084699), (11670,-0.954586), (11671,-0.992155), (11672,-1.235024), (11673,-1.308359), (11674,-1.468087), (11675,-0.788474), (11676,-0.946348), (11677,-0.980197), (11678,-1.155723), (11679,-1.127794), (11680,-1.262443), (11681,-1.358997), (11682,-1.527090), (11683,-0.876738), (11684,-1.068519), (11685,-1.128849), (11686,-1.256065), (11687,-1.003317), (11688,-1.234585), (11689,-1.279116), (11690,-1.451385), (11691,-0.805680), (11692,-0.911069), (11693,-0.976038), (11694,-1.109291), (11695,-1.069753), (11696,-1.215085), (11697,-1.305602), (11698,-1.449074), (11699,-0.788510), (11700,-0.934768), (11701,-0.973727), (11702,-1.119985), (11703,-0.878389), (11704,-1.171434), (11705,-1.227111), (11706,-1.404027), (11707,-0.702586), (11708,-0.877179), (11709,-0.939831), (11710,-1.082370), (11711,-1.110183), (11712,-1.253655), (11713,-1.320484), (11714,-1.473249), (11715,-0.784344), (11716,-0.943614), (11717,-1.039241), (11718,-1.160879), (11719,-0.909533), (11720,-1.134758), (11721,-1.209946), (11722,-1.364101), (11723,-0.643149), (11724,-0.809382), (11725,-0.859029), (11726,-1.008074), (11727,-1.021948), (11728,-1.179822), (11729,-1.248048), (11730,-1.379441), (11731,-0.723053), (11732,-0.852593), (11733,-0.907807), (11734,-1.061961), (11735,-0.833377), (11736,-1.223960), (11737,-1.310764), (11738,-1.472351), (11739,-0.783446), (11740,-0.924595), (11741,-0.983998), (11742,-1.186462), (11743,-1.189653), (11744,-1.328016), (11745,-1.376267), (11746,-1.552719), (11747,-0.877753), (11748,-1.049559), (11749,-1.080158), (11750,-1.222697), (11751,-1.016404), (11752,-1.137585), (11753,-1.203951), (11754,-1.345100), (11755,-0.669201), (11756,-0.846116), (11757,-0.882758), (11758,-1.018797), (11759,-1.038251), (11760,-1.205411), (11761,-1.272240), (11762,-1.433827), (11763,-0.755141), (11764,-0.920911), (11765,-1.041622), (11766,-1.162803), (11767,-0.943505), (11768,-1.112988), (11769,-1.148696), (11770,-1.293558), (11771,-0.607447), (11772,-0.798758), (11773,-0.865124), (11774,-1.026247), (11775,-1.058243), (11776,-1.167344), (11777,-1.236027), (11778,-1.383219), (11779,-0.704070), (11780,-0.868906), (11781,-0.931559), (11782,-1.087573), (11783,-0.858056), (11784,-1.139479), (11785,-1.218857), (11786,-1.400882), (11787,-0.706404), (11788,-0.824329), (11789,-0.885122), (11790,-1.043922), (11791,-1.044791), (11792,-1.188727), (11793,-1.220259), (11794,-1.372553), (11795,-0.716166), (11796,-0.870790), (11797,-0.924613), (11798,-1.078768), (11799,-0.822777), (11800,-0.976931), (11801,-1.139908), (11802,-0.848150), (11803,-1.019956), (11804,-0.655738), (11805,-0.813606), (11806,-0.810298), (11807,-0.958879), (11808,-1.018282), (11809,-1.157108), (11810,-0.889501), (11811,-1.074776), (11812,-0.714271), (11813,-0.905589), (11814,-0.752245), (11815,-0.854378), (11816,-1.114905), (11817,-1.270456), (11818,-1.012135), (11819,-0.779369), (11820,-0.822047), (11821,-0.962732), (11822,-0.953851), (11823,-1.149809), (11824,-1.236613), (11825,-1.328990), (11826,-1.064639), (11827,-0.785880), (11828,-0.826235), (11829,-0.990608), (11830,-0.840521), (11831,-0.933830), (11832,-1.104240), (11833,-1.231457), (11834,-0.959204), (11835,-0.715291), (11836,-0.771438), (11837,-0.903758), (11838,-0.899987), (11839,-1.070403), (11840,-1.152097), (11841,-1.302532), (11842,-1.040505), (11843,-0.827706), (11844,-0.862952), (11845,-1.026399), (11846,-0.890243), (11847,-0.956146), (11848,-1.104264), (11849,-1.273747), (11850,-0.988952), (11851,-0.765941), (11852,-0.797466), (11853,-0.980888), (11854,-0.960855), (11855,-1.121052), (11856,-1.164657), (11857,-1.325317), (11858,-1.046558), (11859,-0.808682), (11860,-0.875981), (11861,-1.007374), (11862,-0.891193), (11863,-0.993326), (11864,-1.007200), (11865,-1.149282), (11866,-0.864957), (11867,-1.000526), (11868,-0.678111), (11869,-0.834589), (11870,-0.820598), (11871,-0.938060), (11872,-1.013718), (11873,-1.144648), (11874,-0.867748), (11875,-0.998215), (11876,-0.686952), (11877,-0.835533), (11878,-0.702628), (11879,-0.827521), (11880,-1.037881), (11881,-1.183212), (11882,-0.884485), (11883,-0.673083), (11884,-0.742699), (11885,-0.908932), (11886,-0.877753), (11887,-1.050486), (11888,-1.093164), (11889,-1.286335), (11890,-0.992717), (11891,-0.727440), (11892,-0.774294), (11893,-0.961429), (11894,-0.821560), (11895,-0.893499), (11896,-1.090853), (11897,-1.244081), (11898,-0.960219), (11899,-0.695862), (11900,-0.759441), (11901,-0.898730), (11902,-0.915860), (11903,-1.116001), (11904,-1.406716), (11905,-1.457290), (11906,-1.201298), (11907,-0.899321), (11908,-1.065085), (11909,-1.154682), (11910,-1.220114), (11911,-1.067704), (11912,-1.330554), (11913,-1.373696), (11914,-1.134423), (11915,-0.833373), (11916,-1.014471), (11917,-1.042747), (11918,-1.247064), (11919,-1.258158), (11920,-1.415562), (11921,-1.413187), (11922,-1.203639), (11923,-0.908631), (11924,-1.057213), (11925,-1.104537), (11926,-1.175079), (11927,-1.037997), (11928,-1.161494), (11929,-1.199995), (11930,-1.368082), (11931,-0.699616), (11932,-0.902548), (11933,-0.949866), (11934,-1.080333), (11935,-1.111395), (11936,-1.263233), (11937,-1.316593), (11938,-1.437767), (11939,-0.801818), (11940,-0.946217), (11941,-1.003296), (11942,-1.162560), (11943,-0.898667), (11944,-1.132720), (11945,-1.311489), (11946,-0.968636), (11947,-1.148808), (11948,-0.866799), (11949,-1.018630), (11950,-1.057132), (11951,-1.208500), (11952,-1.212155), (11953,-1.357487), (11954,-0.991872), (11955,-1.122339), (11956,-0.824538), (11957,-0.975906), (11958,-0.955416), (11959,-1.118394), (11960,-1.234465), (11961,-1.410910), (11962,-1.061094), (11963,-1.201780), (11964,-0.919771), (11965,-1.088791), (11966,-1.163053), (11967,-1.310244), (11968,-1.293461), (11969,-1.421141), (11970,-1.106622), (11971,-1.270069), (11972,-1.005712), (11973,-1.138038), (11974,-1.092458), (11975,-1.275416), (11976,-1.139260), (11977,-1.301781), (11978,-0.954744), (11979,-1.114472), (11980,-0.833396), (11981,-0.975478), (11982,-1.085970), (11983,-1.232228), (11984,-1.243780), (11985,-1.379356), (11986,-1.050904), (11987,-1.184157), (11988,-0.930489), (11989,-1.064669), (11990,-1.054392), (11991,-1.181608), (11992,-1.062178), (11993,-1.214936), (11994,-1.267369), (11995,-1.027633), (11996,-0.751667), (11997,-0.905358), (11998,-0.951286), (11999,-1.104977), (12000,-1.090054), (12001,-1.260470), (12002,-1.294782), (12003,-1.063406), (12004,-0.776757), (12005,-0.953673), (12006,-1.081816), (12007,-1.142146), (12008,-0.986015), (12009,-1.109056), (12010,-1.168452), (12011,-0.946368), (12012,-0.655073), (12013,-0.778107), (12014,-0.804987), (12015,-1.021389), (12016,-1.043628), (12017,-1.201959), (12018,-1.263216), (12019,-1.049027), (12020,-0.748910), (12021,-0.887736), (12022,-0.966644), (12023,-1.020004), (12024,-0.957242), (12025,-1.117896), (12026,-1.135496), (12027,-0.873925), (12028,-0.611428), (12029,-0.782771), (12030,-0.813833), (12031,-0.980066), (12032,-0.897329), (12033,-1.065422), (12034,-1.103454), (12035,-0.846066), (12036,-0.572886), (12037,-0.745156), (12038,-0.829637), (12039,-0.894612), (12040,-0.863434), (12041,-0.999473), (12042,-1.075595), (12043,-0.819597), (12044,-0.565002), (12045,-0.720547), (12046,-0.788309), (12047,-0.978693), (12048,-0.959594), (12049,-1.101669), (12050,-1.157816), (12051,-0.917617), (12052,-0.651406), (12053,-0.801378), (12054,-0.854738), (12055,-0.941542), (12056,-1.090593), (12057,-1.139308), (12058,-1.310650), (12059,-0.634751), (12060,-0.795875), (12061,-0.850625), (12062,-1.003390), (12063,-1.029806), (12064,-1.161206), (12065,-1.246613), (12066,-1.354318), (12067,-0.700254), (12068,-0.833970), (12069,-0.852497), (12070,-1.011761), (12071,-0.782707), (12072,-0.996786), (12073,-1.055719), (12074,-1.205227), (12075,-0.536761), (12076,-0.689062), (12077,-0.750781), (12078,-0.896576), (12079,-0.942968), (12080,-1.062288), (12081,-1.097997), (12082,-1.283272), (12083,-0.638963), (12084,-0.787545), (12085,-0.820003), (12086,-0.974158), (12087,-0.759506), (12088,-1.068800), (12089,-1.116587), (12090,-1.268418), (12091,-0.590203), (12092,-0.750857), (12093,-0.780992), (12094,-0.956518), (12095,-0.949954), (12096,-1.118510), (12097,-1.174194), (12098,-1.332068), (12099,-0.650132), (12100,-0.810323), (12101,-0.874366), (12102,-1.005765), (12103,-0.750701), (12104,-0.983351), (12105,-1.078521), (12106,-1.267972), (12107,-0.556313), (12108,-0.695602), (12109,-0.741530), (12110,-0.891508), (12111,-0.903992), (12112,-1.059543), (12113,-1.102214), (12114,-1.278667), (12115,-0.591622), (12116,-0.748099), (12117,-0.793563), (12118,-0.943078), (12119,-0.697769), (12120,-1.049329), (12121,-1.110122), (12122,-1.262423), (12123,-0.596743), (12124,-0.804316), (12125,-0.886010), (12126,-0.976997), (12127,-0.987621), (12128,-1.145958), (12129,-1.192350), (12130,-1.348827), (12131,-0.643667), (12132,-0.812223), (12133,-0.853042), (12134,-1.019275), (12135,-0.809733), (12136,-1.077223), (12137,-1.155662), (12138,-0.921968), (12139,-0.646929), (12140,-0.808516), (12141,-0.860016), (12142,-1.016494), (12143,-0.990431), (12144,-1.158518), (12145,-1.190977), (12146,-0.987007), (12147,-0.704535), (12148,-0.868445), (12149,-0.872107), (12150,-0.936613), (12151,-0.786525), (12152,-1.197083), (12153,-1.266235), (12154,-1.026036), (12155,-0.770038), (12156,-0.939527), (12157,-0.967803), (12158,-1.127067), (12159,-1.107034), (12160,-0.978781), (12161,-1.033068), (12162,-0.764071), (12163,-0.500178), (12164,-0.661302), (12165,-0.736496), (12166,-0.839092), (12167,-0.694114), (12168,-1.050320), (12169,-0.712576), (12170,-0.872304), (12171,-0.621422), (12172,-0.782082), (12173,-0.848448), (12174,-0.997493), (12175,-0.990935), (12176,-1.141370), (12177,-0.798980), (12178,-0.941989), (12179,-0.648371), (12180,-0.812281), (12181,-0.800614), (12182,-0.938977), (12183,-0.741977), (12184,-0.743778), (12185,-0.940662), (12186,-0.543464), (12187,-0.712020), (12188,-0.422116), (12189,-0.568374), (12190,-0.658898), (12191,-0.811656), (12192,-0.834829), (12193,-1.002452), (12194,-0.625228), (12195,-0.784956), (12196,-0.524781), (12197,-0.663607), (12198,-0.610601), (12199,-0.767078), (12200,-0.896148), (12201,-0.648053), (12202,-0.690731), (12203,-0.840703), (12204,-0.560560), (12205,-0.748158), (12206,-0.805231), (12207,-0.963105), (12208,-0.944469), (12209,-0.715415), (12210,-0.773422), (12211,-0.927113), (12212,-0.670189), (12213,-0.686855), (12214,-0.749038), (12215,-0.897157), (12216,-0.762398), (12217,-0.942100), (12218,-0.626647), (12219,-0.785918), (12220,-0.527597), (12221,-0.656673), (12222,-0.765769), (12223,-0.883230), (12224,-0.904543), (12225,-1.057771), (12226,-0.707015), (12227,-0.841201), (12228,-0.562449), (12229,-0.717530), (12230,-0.675206), (12231,-0.856304), (12232,-0.898512), (12233,-0.607218), (12234,-0.655932), (12235,-0.844463), (12236,-0.552705), (12237,-0.716609), (12238,-0.779725), (12239,-0.930166), (12240,-0.926395), (12241,-0.649496), (12242,-0.709362), (12243,-0.876985), (12244,-0.586617), (12245,-0.681787), (12246,-0.750939), (12247,-0.921812), (12248,-0.833972), (12249,-0.950963), (12250,-0.628548), (12251,-0.774806), (12252,-0.509059), (12253,-0.664610), (12254,-0.741658), (12255,-0.877698), (12256,-0.843269), (12257,-0.985815), (12258,-0.694983), (12259,-0.860284), (12260,-0.586177), (12261,-0.743118), (12262,-0.736561), (12263,-0.876777), (12264,-0.752236), (12265,-0.851583), (12266,-0.477609), (12267,-0.651738), (12268,-0.405496), (12269,-0.545718), (12270,-0.631126), (12271,-0.749983), (12272,-0.735993), (12273,-0.897110), (12274,-0.559367), (12275,-0.711204), (12276,-0.423623), (12277,-0.604258), (12278,-0.594907), (12279,-0.732343), (12280,-0.638454), (12281,-0.772177), (12282,-0.404703), (12283,-0.537492), (12284,-0.257807), (12285,-0.396169), (12286,-0.538714), (12287,-0.708198), (12288,-0.636606), (12289,-0.788907), (12290,-0.443731), (12291,-0.573271), (12292,-0.326102), (12293,-0.470964), (12294,-0.462547), (12295,-0.635749), (12296,-0.670525), (12297,-0.820966), (12298,-0.453492), (12299,-0.603007), (12300,-0.334473), (12301,-0.482122), (12302,-0.569859), (12303,-0.717044), (12304,-0.720235), (12305,-0.865567), (12306,-0.507385), (12307,-0.655504), (12308,-0.395329), (12309,-0.545307), (12310,-0.549426), (12311,-0.694294), (12312,-0.864704), (12313,-0.914815), (12314,-0.680651), (12315,-0.379138), (12316,-0.542121), (12317,-0.580616), (12318,-0.787726), (12319,-0.796960), (12320,-0.967833), (12321,-1.002615), (12322,-0.788427), (12323,-0.501778), (12324,-0.677297), (12325,-0.712543), (12326,-0.755684), (12327,-0.620925), (12328,-0.797377), (12329,-0.856774), (12330,-0.598459), (12331,-0.343395), (12332,-0.507768), (12333,-0.550909), (12334,-0.732934), (12335,-0.733803), (12336,-0.894000), (12337,-0.943178), (12338,-0.640737), (12339,-0.350833), (12340,-0.511956), (12341,-0.584365), (12342,-0.664199), (12343,-0.511325), (12344,-0.772780), (12345,-0.815921), (12346,-0.599873), (12347,-0.312291), (12348,-0.464592), (12349,-0.491935), (12350,-0.666998), (12351,-0.660903), (12352,-0.820167), (12353,-0.892106), (12354,-0.666772), (12355,-0.370831), (12356,-0.512907), (12357,-0.564407), (12358,-0.628920), (12359,-0.503446), (12360,-0.757932), (12361,-0.824761), (12362,-0.599890), (12363,-0.315101), (12364,-0.480401), (12365,-0.505428), (12366,-0.670271), (12367,-0.666493), (12368,-0.818331), (12369,-0.872618), (12370,-0.624053), (12371,-0.354593), (12372,-0.485059), (12373,-0.550962), (12374,-0.631723), (12375,-0.468630), (12376,-0.811374), (12377,-0.866124), (12378,-0.638930), (12379,-0.347172), (12380,-0.497144), (12381,-0.555150), (12382,-0.724170), (12383,-0.729685), (12384,-0.889418), (12385,-0.949742), (12386,-0.705359), (12387,-0.435899), (12388,-0.611888), (12389,-0.641091), (12390,-0.722322), (12391,-0.553186), (12392,-0.918691), (12393,-0.597202), (12394,-0.730455), (12395,-0.462385), (12396,-0.626295), (12397,-0.750256), (12398,-0.893265), (12399,-0.903426), (12400,-1.049221), (12401,-0.688253), (12402,-0.844730), (12403,-0.566904), (12404,-0.698304), (12405,-0.674558), (12406,-0.808738), (12407,-0.663296), (12408,-0.822560), (12409,-0.907041), (12410,-0.687280), (12411,-0.382510), (12412,-0.547353), (12413,-0.579812), (12414,-0.750685), (12415,-0.698142), (12416,-0.869021), (12417,-1.034784), (12418,-0.483837), (12419,-0.599438), (12420,-0.676023), (12421,-0.821818), (12422,-0.478038), (12423,-0.642875), (12424,-0.822114), (12425,-0.851323), (12426,-0.613440), (12427,-0.613389), (12428,-0.771256), (12429,-0.821367), (12430,-0.975985), (12431,-0.713024), (12432,-0.854173), (12433,-0.891278), (12434,-0.646896), (12435,-0.507490), (12436,-0.669541), (12437,-0.714542), (12438,-0.777658), (12439,-0.516557), (12440,-0.806809), (12441,-0.873175), (12442,-0.614854), (12443,-0.574389), (12444,-0.774530), (12445,-0.820457), (12446,-0.996910), (12447,-0.714438), (12448,-0.874171), (12449,-0.943323), (12450,-0.697082), (12451,-0.526092), (12452,-0.672351), (12453,-0.752649), (12454,-0.831093), (12455,-0.550481), (12456,-0.955002), (12457,-0.628868), (12458,-0.806716), (12459,-0.768569), (12460,-0.916223), (12461,-1.016960), (12462,-1.141390), (12463,-0.866351), (12464,-1.048376), (12465,-0.682298), (12466,-0.811831), (12467,-0.668250), (12468,-0.829373), (12469,-0.808877), (12470,-0.949563), (12471,-0.692175), (12472,-0.908107), (12473,-0.926164), (12474,-0.709189), (12475,-0.699845), (12476,-0.869792), (12477,-0.964028), (12478,-1.141870), (12479,-0.858935), (12480,-1.015882), (12481,-1.045548), (12482,-0.816964), (12483,-0.666407), (12484,-0.810349), (12485,-0.899006), (12486,-0.935184), (12487,-0.636457), (12488,-0.833341), (12489,-0.878342), (12490,-0.661367), (12491,-0.645981), (12492,-0.795026), (12493,-0.857678), (12494,-1.038777), (12495,-0.748872), (12496,-0.900704), (12497,-0.949887), (12498,-0.692036), (12499,-0.515468), (12500,-0.687274), (12501,-0.741098), (12502,-0.810250), (12503,-0.551472), (12504,-0.853340), (12505,-0.935961), (12506,-0.694365), (12507,-0.671082), (12508,-0.819664), (12509,-0.828435), (12510,-1.021606), (12511,-0.756322), (12512,-0.912336), (12513,-0.981958), (12514,-0.716211), (12515,-0.554508), (12516,-0.707736), (12517,-0.784321), (12518,-0.846967), (12519,-0.581683), (12520,-0.705650), (12521,-0.755291), (12522,-0.519274), (12523,-0.525716), (12524,-0.662225), (12525,-0.768071), (12526,-0.940340), (12527,-0.671343), (12528,-0.841753), (12529,-0.865853), (12530,-0.618684), (12531,-0.493217), (12532,-0.652945), (12533,-0.680294), (12534,-0.753159), (12535,-0.450255), (12536,-0.762799), (12537,-0.824988), (12538,-0.581533), (12539,-0.581481), (12540,-0.765823), (12541,-0.818257), (12542,-0.984026), (12543,-0.714097), (12544,-0.830161), (12545,-0.830573), (12546,-0.595483), (12547,-0.414268), (12548,-0.562850), (12549,-0.625503), (12550,-0.684436), (12551,-0.414506), (12552,-0.732165), (12553,-0.785989), (12554,-0.546716), (12555,-0.527617), (12556,-0.689667), (12557,-0.793659), (12558,-0.973361), (12559,-0.671384), (12560,-0.830185), (12561,-0.884008), (12562,-0.647986), (12563,-0.472820), (12564,-0.636260), (12565,-0.703559), (12566,-0.789893), (12567,-0.515324), (12568,-0.674588), (12569,-0.826419), (12570,-0.806393), (12571,-0.558297), (12572,-0.627449), (12573,-0.795073), (12574,-0.505638), (12575,-0.695096), (12576,-0.692714), (12577,-0.842223), (12578,-0.687026), (12579,-0.451009), (12580,-0.498790), (12581,-0.604642), (12582,-0.327280), (12583,-0.383426), (12584,-0.633265), (12585,-0.800895), (12586,-0.409733), (12587,-0.557851), (12588,-0.637686), (12589,-0.802059), (12590,-0.545605), (12591,-0.641231), (12592,-0.699238), (12593,-0.847356), (12594,-0.341461), (12595,-0.511414), (12596,-0.551762), (12597,-0.719855), (12598,-0.345418), (12599,-0.510718), (12600,-0.787965), (12601,-0.929577), (12602,-0.508227), (12603,-0.681424), (12604,-0.746399), (12605,-0.897304), (12606,-0.649202), (12607,-0.808473), (12608,-0.860900), (12609,-1.011805), (12610,-0.431596), (12611,-0.584824), (12612,-0.651653), (12613,-0.772827), (12614,-0.413719), (12615,-0.560904), (12616,-0.706236), (12617,-0.832983), (12618,-0.442754), (12619,-0.599695), (12620,-0.661414), (12621,-0.822538), (12622,-0.567473), (12623,-0.742529), (12624,-0.792177), (12625,-0.927289), (12626,-0.365190), (12627,-0.549538), (12628,-0.619160), (12629,-0.759839), (12630,-0.389585), (12631,-0.560928), (12632,-0.609642), (12633,-0.782375), (12634,-0.717289), (12635,-0.525862), (12636,-0.608020), (12637,-0.722694), (12638,-0.443472), (12639,-0.642685), (12640,-0.716484), (12641,-0.904545), (12642,-0.730770), (12643,-0.493820), (12644,-0.536035), (12645,-0.687866), (12646,-0.389602), (12647,-0.488021), (12648,-0.846087), (12649,-0.472577), (12650,-0.622085), (12651,-0.635039), (12652,-0.783620), (12653,-0.827225), (12654,-0.969301), (12655,-0.696121), (12656,-0.837270), (12657,-0.491167), (12658,-0.667619), (12659,-0.526818), (12660,-0.683295), (12661,-0.648403), (12662,-0.832288), (12663,-0.543780), (12664,-0.722555), (12665,-0.888782), (12666,-0.473469), (12667,-0.668036), (12668,-0.714427), (12669,-0.856509), (12670,-0.576360), (12671,-0.706364), (12672,-0.899071), (12673,-0.960791), (12674,-0.698294), (12675,-0.593728), (12676,-0.725585), (12677,-0.759440), (12678,-0.850421), (12679,-0.568882), (12680,-0.788070), (12681,-0.830741), (12682,-0.599371), (12683,-0.585844), (12684,-0.749285), (12685,-0.810541), (12686,-0.966555), (12687,-0.678980), (12688,-0.861005), (12689,-0.900890), (12690,-0.654655), (12691,-0.541724), (12692,-0.676836), (12693,-0.742275), (12694,-0.790526), (12695,-0.498762), (12696,-0.767186), (12697,-0.926450), (12698,-0.596138), (12699,-0.761902), (12700,-0.754881), (12701,-0.883024), (12702,-0.947067), (12703,-1.116087), (12704,-0.811787), (12705,-0.978947), (12706,-0.667677), (12707,-0.797217), (12708,-0.636910), (12709,-0.798034), (12710,-0.789147), (12711,-0.936802), (12712,-0.711931), (12713,-0.886060), (12714,-0.540884), (12715,-0.693179), (12716,-0.670829), (12717,-0.829166), (12718,-0.914574), (12719,-1.088240), (12720,-0.797408), (12721,-0.925552), (12722,-0.589198), (12723,-0.722451), (12724,-0.590478), (12725,-0.730237), (12726,-0.691163), (12727,-0.837421), (12728,-0.729600), (12729,-0.890724), (12730,-0.579454), (12731,-0.706671), (12732,-0.672706), (12733,-0.851018), (12734,-0.927603), (12735,-1.048777), (12736,-0.765842), (12737,-0.939508), (12738,-0.598508), (12739,-0.727121), (12740,-0.602111), (12741,-0.754876), (12742,-0.735776), (12743,-0.884357), (12744,-0.675742), (12745,-0.798776), (12746,-0.464282), (12747,-0.612863), (12748,-0.629994), (12749,-0.774856), (12750,-0.877921), (12751,-0.980054), (12752,-0.718947), (12753,-0.872638), (12754,-0.534431), (12755,-0.688585), (12756,-0.544534), (12757,-0.701944), (12758,-0.644291), (12759,-0.814701), (12760,-0.778876), (12761,-0.938140), (12762,-0.592037), (12763,-0.731796), (12764,-0.729878), (12765,-0.895648), (12766,-1.005677), (12767,-1.164014), (12768,-0.870859), (12769,-1.036629), (12770,-0.664046), (12771,-0.833992), (12772,-0.687617), (12773,-0.825517), (12774,-0.798521), (12775,-0.952675), (12776,-0.699007), (12777,-0.832723), (12778,-0.513095), (12779,-0.649597), (12780,-0.622138), (12781,-0.756781), (12782,-0.860774), (12783,-0.999600), (12784,-0.712488), (12785,-0.868032), (12786,-0.545617), (12787,-0.703954), (12788,-0.568732), (12789,-0.762829), (12790,-0.719578), (12791,-0.892775), (12792,-0.665581), (12793,-0.812772), (12794,-0.443438), (12795,-0.603635), (12796,-0.591035), (12797,-0.760518), (12798,-0.844999), (12799,-1.013092), (12800,-0.744095), (12801,-0.894067), (12802,-0.517770), (12803,-0.672851), (12804,-0.545525), (12805,-0.703862), (12806,-0.634594), (12807,-0.761810), (12808,-0.659098), (12809,-0.812789), (12810,-0.457394), (12811,-0.649175), (12812,-0.639361), (12813,-0.808851), (12814,-0.879856), (12815,-1.021005), (12816,-0.741789), (12817,-0.888048), (12818,-0.557273), (12819,-0.709568), (12820,-0.572486), (12821,-0.717818), (12822,-0.677816), (12823,-0.823605), (12824,-0.639147), (12825,-0.670673), (12826,-0.833656), (12827,-0.440171), (12828,-0.605941), (12829,-0.655582), (12830,-0.845973), (12831,-0.558391), (12832,-0.704186), (12833,-0.787271), (12834,-0.907518), (12835,-0.379795), (12836,-0.520481), (12837,-0.567805), (12838,-0.717783), (12839,-0.341480), (12840,-0.759933), (12841,-0.823049), (12842,-0.581923), (12843,-0.568860), (12844,-0.701180), (12845,-0.769869), (12846,-0.971868), (12847,-0.681037), (12848,-0.824509), (12849,-0.878803), (12850,-0.652535), (12851,-0.470394), (12852,-0.636627), (12853,-0.689061), (12854,-0.787011), (12855,-0.487820), (12856,-0.765993), (12857,-0.814244), (12858,-0.589836), (12859,-0.570273), (12860,-0.777376), (12861,-0.834456), (12862,-1.013232), (12863,-0.723790), (12864,-0.894206), (12865,-0.936415), (12866,-0.687392), (12867,-0.537305), (12868,-0.680307), (12869,-0.767111), (12870,-0.851129), (12871,-0.569126), (12872,-0.808283), (12873,-0.840278), (12874,-0.596823), (12875,-0.592588), (12876,-0.744883), (12877,-0.768056), (12878,-0.927320), (12879,-0.636025), (12880,-0.808295), (12881,-0.845393), (12882,-0.601017), (12883,-0.457893), (12884,-0.602761), (12885,-0.662621), (12886,-0.750821), (12887,-0.463703), (12888,-0.605322), (12889,-0.652176), (12890,-0.803081), (12891,-0.395663), (12892,-0.531703), (12893,-0.610147), (12894,-0.754546), (12895,-0.496232), (12896,-0.683830), (12897,-0.720935), (12898,-0.866260), (12899,-0.338537), (12900,-0.490375), (12901,-0.556741), (12902,-0.700213), (12903,-0.326703), (12904,-0.726108), (12905,-0.774359), (12906,-0.552738), (12907,-0.518773), (12908,-0.666891), (12909,-0.734653), (12910,-0.905989), (12911,-0.610055), (12912,-0.782788), (12913,-0.832898), (12914,-0.575047), (12915,-0.429136), (12916,-0.609765), (12917,-0.637114), (12918,-0.719742), (12919,-0.441452), (12920,-0.745173), (12921,-0.817112), (12922,-0.585272), (12923,-0.555026), (12924,-0.722186), (12925,-0.752322), (12926,-0.934810), (12927,-0.655131), (12928,-1.052677), (12929,-1.082813), (12930,-0.863051), (12931,-0.718073), (12932,-0.870368), (12933,-0.937197), (12934,-0.974302), (12935,-0.751291), (12936,-0.828803), (12937,-0.966702), (12938,-0.624775), (12939,-0.770107), (12940,-0.744501), (12941,-0.906552), (12942,-0.989642), (12943,-1.138224), (12944,-0.872477), (12945,-1.060538), (12946,-0.720935), (12947,-0.820744), (12948,-0.642786), (12949,-0.798800), (12950,-0.756939), (12951,-0.903661), (12952,-0.855764), (12953,-0.994126), (12954,-0.649877), (12955,-0.809610), (12956,-0.815588), (12957,-0.949774), (12958,-1.006385), (12959,-1.159612), (12960,-0.892469), (12961,-1.065202), (12962,-0.722812), (12963,-0.861174), (12964,-0.744530), (12965,-0.882893), (12966,-0.856824), (12967,-1.000296), (12968,-0.780534), (12969,-0.897069), (12970,-0.554679), (12971,-0.722766), (12972,-0.709239), (12973,-0.863393), (12974,-0.933015), (12975,-1.079737), (12976,-0.802844), (12977,-0.951426), (12978,-0.620181), (12979,-0.752508), (12980,-0.607530), (12981,-0.773293), (12982,-0.742578), (12983,-0.906025), (12984,-0.863237), (12985,-1.022038), (12986,-0.674075), (12987,-0.800822), (12988,-0.827708), (12989,-0.976290), (12990,-1.055661), (12991,-1.187987), (12992,-0.918984), (12993,-1.082894), (12994,-0.752120), (12995,-0.941577), (12996,-0.803099), (12997,-0.911268), (12998,-0.924221), (12999,-1.058864), (13000,-0.730876), (13001,-0.894323), (13002,-0.551933), (13003,-0.708411), (13004,-0.673513), (13005,-0.837423), (13006,-0.932592), (13007,-1.042621), (13008,-0.756899), (13009,-0.947747), (13010,-0.645770), (13011,-0.798065), (13012,-0.634045), (13013,-0.777517), (13014,-0.750051), (13015,-0.945552), (13016,-0.894398), (13017,-1.056449), (13018,-0.710809), (13019,-0.870073), (13020,-0.839358), (13021,-0.987013), (13022,-1.063134), (13023,-1.220539), (13024,-0.939926), (13025,-1.057387), (13026,-0.706175), (13027,-0.869152), (13028,-0.700486), (13029,-0.876475), (13030,-0.835077), (13031,-0.976226), (13032,-0.672389), (13033,-0.856274), (13034,-0.521317), (13035,-0.672685), (13036,-0.678663), (13037,-0.855579), (13038,-0.906153), (13039,-1.053807), (13040,-0.757403), (13041,-0.925490), (13042,-0.595179), (13043,-0.765125), (13044,-0.616897), (13045,-0.799386), (13046,-0.755202), (13047,-0.892174), (13048,-0.502402), (13049,-0.683964), (13050,-0.728502), (13051,-0.485046), (13052,-0.455264), (13053,-0.632643), (13054,-0.692509), (13055,-0.890326), (13056,-0.546540), (13057,-0.693731), (13058,-0.776352), (13059,-0.544512), (13060,-0.378633), (13061,-0.494234), (13062,-0.551777), (13063,-0.644154), (13064,-0.494066), (13065,-0.673305), (13066,-0.713654), (13067,-0.486460), (13068,-0.458537), (13069,-0.625234), (13070,-0.669302), (13071,-0.852254), (13072,-0.571648), (13073,-0.722546), (13074,-0.778229), (13075,-0.538030), (13076,-0.387016), (13077,-0.566254), (13078,-0.605676), (13079,-0.683657), (13080,-0.641327), (13081,-0.691901), (13082,-0.857671), (13083,-0.457686), (13084,-0.621596), (13085,-0.690285), (13086,-0.836074), (13087,-0.586588), (13088,-0.738883), (13089,-0.818254), (13090,-0.959403), (13091,-0.424248), (13092,-0.551001), (13093,-0.602038), (13094,-0.750156), (13095,-0.366427), (13096,-0.774198), (13097,-0.806650), (13098,-0.554842), (13099,-0.545492), (13100,-0.715908), (13101,-0.763695), (13102,-0.922959), (13103,-0.631195), (13104,-0.783032), (13105,-0.851252), (13106,-0.617095), (13107,-0.468860), (13108,-0.627198), (13109,-0.692637), (13110,-0.786867), (13111,-0.516944), (13112,-0.668312), (13113,-0.726318), (13114,-0.880936), (13115,-0.497206), (13116,-0.598875), (13117,-0.668491), (13118,-0.813360), (13119,-0.562008), (13120,-0.704553), (13121,-0.774169), (13122,-0.963163), (13123,-0.415002), (13124,-0.574730), (13125,-0.623444), (13126,-0.788287), (13127,-0.444037), (13128,-0.639995), (13129,-0.706830), (13130,-0.854479), (13131,-0.473072), (13132,-0.648128), (13133,-0.693593), (13134,-0.808731), (13135,-0.540660), (13136,-0.706894), (13137,-0.778832), (13138,-0.903263), (13139,-0.374143), (13140,-0.506933), (13141,-0.535679), (13142,-0.680077), (13143,-0.318646), (13144,-0.594033), (13145,-0.664111), (13146,-0.821522), (13147,-0.433610), (13148,-0.578015), (13149,-0.641124), (13150,-0.825473), (13151,-0.565299), (13152,-0.718990), (13153,-0.763064), (13154,-0.911176), (13155,-0.374630), (13156,-0.520425), (13157,-0.575176), (13158,-0.710288), (13159,-0.351180), (13160,-0.599629), (13161,-0.759356), (13162,-0.429045), (13163,-0.592022), (13164,-0.613799), (13165,-0.751698), (13166,-0.812021), (13167,-0.982901), (13168,-0.713440), (13169,-0.878277), (13170,-0.547496), (13171,-0.685859), (13172,-0.548777), (13173,-0.708510), (13174,-0.658284), (13175,-0.809188), (13176,-0.889029), (13177,-0.972577), (13178,-0.699861), (13179,-0.686804), (13180,-0.818660), (13181,-0.849259), (13182,-1.034071), (13183,-0.778080), (13184,-0.770589), (13185,-0.924280), (13186,-0.947447), (13187,-0.704461), (13188,-0.553446), (13189,-0.711777), (13190,-0.793941), (13191,-0.855661), (13192,-0.680026), (13193,-0.833717), (13194,-0.859670), (13195,-0.648268), (13196,-0.618949), (13197,-0.780999), (13198,-0.823214), (13199,-0.985264), (13200,-0.711158), (13201,-0.908042), (13202,-0.944220), (13203,-0.674754), (13204,-0.535349), (13205,-0.683930), (13206,-0.738217), (13207,-0.812016), (13208,-0.649386), (13209,-0.798431), (13210,-0.835072), (13211,-0.616701), (13212,-0.605961), (13213,-0.768017), (13214,-0.841810), (13215,-0.987605), (13216,-0.704206), (13217,-0.889018), (13218,-0.992083), (13219,-0.739342), (13220,-0.592504), (13221,-0.748054), (13222,-0.803268), (13223,-0.855702), (13224,-0.823597), (13225,-0.941984), (13226,-0.617246), (13227,-0.780693), (13228,-0.762520), (13229,-0.897626), (13230,-0.956096), (13231,-1.121866), (13232,-0.851473), (13233,-1.013993), (13234,-0.699937), (13235,-0.857341), (13236,-0.758812), (13237,-0.909253), (13238,-0.841375), (13239,-0.997389), (13240,-0.805035), (13241,-0.941075), (13242,-0.965638), (13243,-0.718006), (13244,-0.694260), (13245,-0.821470), (13246,-0.919426), (13247,-1.063362), (13248,-0.788786), (13249,-0.944800), (13250,-0.965180), (13251,-0.763534), (13252,-0.600904), (13253,-0.758308), (13254,-0.824674), (13255,-0.897082), (13256,-0.655486), (13257,-0.790136), (13258,-0.840710), (13259,-0.615369), (13260,-0.613921), (13261,-0.758783), (13262,-0.810753), (13263,-0.960262), (13264,-0.699161), (13265,-0.860284), (13266,-0.937796), (13267,-0.706889), (13268,-0.564691), (13269,-0.747649), (13270,-0.779175), (13271,-0.839505), (13272,-0.742365), (13273,-0.866796), (13274,-0.941521), (13275,-0.715260), (13276,-0.705910), (13277,-0.864247), (13278,-0.897169), (13279,-1.064792), (13280,-0.786503), (13281,-0.925329), (13282,-0.983799), (13283,-0.708303), (13284,-0.564251), (13285,-0.727228), (13286,-0.780125), (13287,-0.834882), (13288,-0.856189), (13289,-0.591368), (13290,-0.751565), (13291,-0.445869), (13292,-0.574945), (13293,-0.566991), (13294,-0.704890), (13295,-0.777293), (13296,-0.914728), (13297,-0.635969), (13298,-0.832860), (13299,-0.489080), (13300,-0.648344), (13301,-0.482928), (13302,-0.635686), (13303,-0.614263), (13304,-0.598883), (13305,-0.707978), (13306,-0.783636), (13307,-0.553186), (13308,-0.508075), (13309,-0.639469), (13310,-0.700725), (13311,-0.898079), (13312,-0.617003), (13313,-0.808784), (13314,-0.857035), (13315,-0.613585), (13316,-0.485326), (13317,-0.616719), (13318,-0.669153), (13319,-0.754097), (13320,-0.951914), (13321,-0.664339), (13322,-0.817560), (13323,-0.467744), (13324,-0.624685), (13325,-0.625554), (13326,-0.768562), (13327,-0.828429), (13328,-0.950529), (13329,-0.688502), (13330,-0.860308), (13331,-0.510949), (13332,-0.655354), (13333,-0.519198), (13334,-0.627367), (13335,-0.622669), (13336,-0.671383), (13337,-0.705696), (13338,-0.863106), (13339,-0.427348), (13340,-0.593582), (13341,-0.634870), (13342,-0.782518), (13343,-0.544178), (13344,-0.702516), (13345,-0.761449), (13346,-0.930932), (13347,-0.422251), (13348,-0.550394), (13349,-0.581926), (13350,-0.775097), (13351,-0.437353), (13352,-0.545522), (13353,-0.703859), (13354,-0.734459), (13355,-0.503082), (13356,-0.481659), (13357,-0.628387), (13358,-0.675242), (13359,-0.859590), (13360,-0.580374), (13361,-0.710371), (13362,-0.745153), (13363,-0.529105), (13364,-0.392955), (13365,-0.561042), (13366,-0.605580), (13367,-0.707712), (13368,-0.722519), (13369,-0.771697), (13370,-0.916096), (13371,-0.531903), (13372,-0.670265), (13373,-0.700864), (13374,-0.855489), (13375,-0.615283), (13376,-0.777803), (13377,-0.819548), (13378,-0.977885), (13379,-0.430651), (13380,-0.594098), (13381,-0.643281), (13382,-0.818337), (13383,-0.424852), (13384,-0.598055), (13385,-0.793549), (13386,-0.829721), (13387,-0.619715), (13388,-0.605255), (13389,-0.758946), (13390,-0.790015), (13391,-0.952065), (13392,-0.661697), (13393,-0.780085), (13394,-0.889187), (13395,-0.636445), (13396,-0.481248), (13397,-0.646085), (13398,-0.698982), (13399,-0.732368), (13400,-0.652417), (13401,-0.714606), (13402,-0.881766), (13403,-0.479458), (13404,-0.617821), (13405,-0.666998), (13406,-0.835091), (13407,-0.563302), (13408,-0.687269), (13409,-0.746202), (13410,-0.963061), (13411,-0.380529), (13412,-0.530971), (13413,-0.605232), (13414,-0.744058), (13415,-0.389126), (13416,-0.651977), (13417,-0.833533), (13418,-0.475351), (13419,-0.625329), (13420,-0.601119), (13421,-0.771992), (13422,-0.870412), (13423,-1.003201), (13424,-0.742094), (13425,-0.894395), (13426,-0.529707), (13427,-0.667607), (13428,-0.513336), (13429,-0.676783), (13430,-0.652110), (13431,-0.796972), (13432,-0.572102), (13433,-0.738798), (13434,-0.797268), (13435,-0.559392), (13436,-0.523567), (13437,-0.680508), (13438,-0.711570), (13439,-0.913107), (13440,-0.779738), (13441,-0.924143), (13442,-0.965424), (13443,-0.760528), (13444,-0.611831), (13445,-0.745084), (13446,-0.792408), (13447,-0.888961), (13448,-0.716582), (13449,-0.874450), (13450,-0.924097), (13451,-0.683897), (13452,-0.619275), (13453,-0.798044), (13454,-0.848618), (13455,-1.051545), (13456,-0.794163), (13457,-0.924160), (13458,-0.977520), (13459,-0.718743), (13460,-0.577014), (13461,-0.735815), (13462,-0.782669), (13463,-0.845322), (13464,-0.652035), (13465,-0.821055), (13466,-0.909249), (13467,-0.674159), (13468,-0.710337), (13469,-0.865418), (13470,-0.883939), (13471,-1.055281), (13472,-0.775139), (13473,-0.940439), (13474,-0.966862), (13475,-0.745241), (13476,-0.601189), (13477,-0.757203), (13478,-0.824959), (13479,-0.881106), (13480,-1.172291), (13481,-0.910257), (13482,-0.654266), (13483,-0.704370), (13484,-0.864567), (13485,-0.851503), (13486,-1.005658), (13487,-1.042299), (13488,-1.220142), (13489,-0.933493), (13490,-0.701653), (13491,-0.729003), (13492,-0.917064), (13493,-0.768836), (13494,-0.840311), (13495,-0.911787), (13496,-1.118426), (13497,-0.824809), (13498,-0.979433), (13499,-0.607312), (13500,-0.759144), (13501,-0.758622), (13502,-0.920216), (13503,-0.987508), (13504,-1.154668), (13505,-0.836436), (13506,-0.980835), (13507,-0.647267), (13508,-0.798642), (13509,-0.668059), (13510,-0.813854), (13511,-0.776170), (13512,-0.962378), (13513,-0.673406), (13514,-0.840566), (13515,-0.501432), (13516,-0.658837), (13517,-0.641590), (13518,-0.781812), (13519,-0.861184), (13520,-0.965639), (13521,-0.726830), (13522,-0.887490), (13523,-0.565538), (13524,-0.686719), (13525,-0.558923), (13526,-0.694962), (13527,-0.669357), (13528,-0.998631), (13529,-0.725915), (13530,-0.886575), (13531,-0.531180), (13532,-0.686261), (13533,-0.684350), (13534,-0.838041), (13535,-0.938314), (13536,-1.087358), (13537,-0.829507), (13538,-0.971120), (13539,-0.657997), (13540,-0.830730), (13541,-0.692721), (13542,-0.848265), (13543,-0.836598), (13544,-0.961022), (13545,-0.689702), (13546,-0.855472), (13547,-0.520978), (13548,-0.655158), (13549,-0.640241), (13550,-0.800432), (13551,-0.892808), (13552,-1.045573), (13553,-0.731054), (13554,-0.848051), (13555,-0.494516), (13556,-0.666785), (13557,-0.525520), (13558,-0.649017), (13559,-0.609943), (13560,-0.915523), (13561,-0.650240), (13562,-0.813686), (13563,-0.474546), (13564,-0.653322), (13565,-0.635149), (13566,-0.778621), (13567,-0.837090), (13568,-1.071607), (13569,-0.786812), (13570,-0.960015), (13571,-0.616692), (13572,-0.770852), (13573,-0.610076), (13574,-0.752621), (13575,-0.726552), (13576,-1.065113), (13577,-0.767313), (13578,-0.920077), (13579,-0.607417), (13580,-0.734165), (13581,-0.694627), (13582,-0.835776), (13583,-0.907714), (13584,-1.072088), (13585,-0.794268), (13586,-0.927521), (13587,-0.594417), (13588,-0.758328), (13589,-0.612423), (13590,-0.746602), (13591,-0.751191), (13592,-0.558367), (13593,-0.677688), (13594,-0.755669), (13595,-0.899141), (13596,-0.491717), (13597,-0.637512), (13598,-0.708988), (13599,-0.859429), (13600,-0.602041), (13601,-0.746440), (13602,-0.842073), (13603,-0.980436), (13604,-0.436921), (13605,-0.559491), (13606,-0.633753), (13607,-0.793944), (13608,-0.593694), (13609,-0.765500), (13610,-0.833256), (13611,-0.614421), (13612,-0.586029), (13613,-0.730434), (13614,-0.810269), (13615,-0.990904), (13616,-0.698213), (13617,-0.822173), (13618,-0.902014), (13619,-0.665528), (13620,-0.547951), (13621,-0.656126), (13622,-0.687652), (13623,-0.751695), (13624,-0.683359), (13625,-0.843087), (13626,-0.901093), (13627,-0.666003), (13628,-0.648757), (13629,-0.813130), (13630,-0.864174), (13631,-1.054095), (13632,-0.764654), (13633,-0.960148), (13634,-0.995863), (13635,-0.749158), (13636,-0.582345), (13637,-0.748578), (13638,-0.765708), (13639,-0.850189), (13640,-0.704748), (13641,-0.865402), (13642,-0.912726), (13643,-0.679959), (13644,-0.645061), (13645,-0.791789), (13646,-0.827035), (13647,-0.988152), (13648,-0.721015), (13649,-0.896071), (13650,-0.936426), (13651,-0.695293), (13652,-0.557284), (13653,-0.710975), (13654,-0.751330), (13655,-0.820946), (13656,-0.463227), (13657,-0.627601), (13658,-0.687467), (13659,-0.853700), (13660,-0.440704), (13661,-0.617156), (13662,-0.669589), (13663,-0.834890), (13664,-0.566820), (13665,-0.695896), (13666,-0.740891), (13667,-0.881576), (13668,-0.369652), (13669,-0.507081), (13670,-0.569734), (13671,-0.718779), (13672,-0.690850), (13673,-0.855693), (13674,-0.519339), (13675,-0.679067), (13676,-0.665540), (13677,-0.837809), (13678,-0.893029), (13679,-1.027679), (13680,-0.739634), (13681,-0.877996), (13682,-0.580196), (13683,-0.731101), (13684,-0.590305), (13685,-0.768148), (13686,-0.713744), (13687,-0.848394), (13688,-0.628163), (13689,-0.789750), (13690,-0.836611), (13691,-0.595478), (13692,-0.566623), (13693,-0.702662), (13694,-0.752773), (13695,-0.930152), (13696,-0.701098), (13697,-0.870118), (13698,-0.952282), (13699,-0.699071), (13700,-0.578713), (13701,-0.738904), (13702,-0.801557), (13703,-0.885111), (13704,-0.665343), (13705,-0.832509), (13706,-0.877504), (13707,-0.625696), (13708,-0.636783), (13709,-0.785365), (13710,-0.849408), (13711,-1.032829), (13712,-0.753144), (13713,-0.891043), (13714,-0.953695), (13715,-0.735324), (13716,-0.593132), (13717,-0.692942), (13718,-0.762557), (13719,-0.817314), (13720,-0.965426), (13721,-0.705722), (13722,-0.851047), (13723,-0.524455), (13724,-0.671177), (13725,-0.673906), (13726,-0.845712), (13727,-0.922297), (13728,-1.092243), (13729,-0.803741), (13730,-0.955572), (13731,-0.621078), (13732,-0.752472), (13733,-0.619572), (13734,-0.763971), (13735,-0.686807), (13736,-1.162861), (13737,-0.909187), (13738,-0.662951), (13739,-0.689367), (13740,-0.836096), (13741,-0.810490), (13742,-1.009697), (13743,-1.064917), (13744,-1.214425), (13745,-0.912912), (13746,-0.699656), (13747,-0.760913), (13748,-0.928072), (13749,-0.747791), (13750,-0.793719), (13751,-0.858231), (13752,-1.059298), (13753,-0.797727), (13754,-0.908689), (13755,-0.568159), (13756,-0.742751), (13757,-0.744553), (13758,-0.913573), (13759,-0.970646), (13760,-1.102039), (13761,-0.858127), (13762,-0.984874), (13763,-0.655026), (13764,-0.837978), (13765,-0.693933), (13766,-0.816034), (13767,-0.767673), (13768,-0.997538), (13769,-0.700207), (13770,-0.878519), (13771,-0.519404), (13772,-0.652657), (13773,-0.624265), (13774,-0.844843), (13775,-0.924684), (13776,-1.073266), (13777,-0.755490), (13778,-0.910578), (13779,-0.581193), (13780,-0.723269), (13781,-0.603375), (13782,-0.755206), (13783,-0.702200), (13784,-1.031931), (13785,-0.728558), (13786,-0.894791), (13787,-0.535219), (13788,-0.695873), (13789,-0.688852), (13790,-0.821642), (13791,-0.898227), (13792,-1.035193), (13793,-0.779665), (13794,-0.940325), (13795,-0.569601), (13796,-0.715860), (13797,-0.570882), (13798,-0.727823), (13799,-0.722192), (13800,-0.876346), (13801,-0.614782), (13802,-0.751285), (13803,-0.413078), (13804,-0.574665), (13805,-0.563924), (13806,-0.721328), (13807,-0.806273), (13808,-0.954391), (13809,-0.651487), (13810,-0.822830), (13811,-0.479507), (13812,-0.640167), (13813,-0.493329), (13814,-0.647020), (13815,-0.631170), (13816,-0.937214), (13817,-0.636170), (13818,-0.771277), (13819,-0.413095), (13820,-0.562609), (13821,-0.590422), (13822,-0.757582), (13823,-0.867610), (13824,-0.918184), (13825,-0.640822), (13826,-0.822384), (13827,-0.513437), (13828,-0.640184), (13829,-0.502639), (13830,-0.646111), (13831,-0.613079), (13832,-0.948384), (13833,-0.674741), (13834,-0.822395), (13835,-0.455848), (13836,-0.605363), (13837,-0.639211), (13838,-0.814731), (13839,-0.889925), (13840,-1.048263), (13841,-0.785302), (13842,-0.888361), (13843,-0.556654), (13844,-0.709418), (13845,-0.579299), (13846,-0.734386), (13847,-0.722719), (13848,-0.648341), (13849,-0.815501), (13850,-0.846101), (13851,-0.601725), (13852,-0.575656), (13853,-0.707976), (13854,-0.746471), (13855,-0.951720), (13856,-0.663218), (13857,-0.879614), (13858,-0.944583), (13859,-0.676513), (13860,-0.504134), (13861,-0.671294), (13862,-0.749269), (13863,-0.775228), (13864,-0.521554), (13865,-0.672458), (13866,-0.732324), (13867,-0.474937), (13868,-0.482775), (13869,-0.649935), (13870,-0.700045), (13871,-0.838871), (13872,-0.530858), (13873,-0.687335), (13874,-0.744872), (13875,-0.509319), (13876,-0.364341), (13877,-0.517099), (13878,-0.570459), (13879,-0.661909), (13880,-0.607043), (13881,-0.779775), (13882,-0.825703), (13883,-0.567852), (13884,-0.571514), (13885,-0.724278), (13886,-0.753944), (13887,-0.958267), (13888,-0.674405), (13889,-0.844351), (13890,-0.892602), (13891,-0.646830), (13892,-0.510674), (13893,-0.646714), (13894,-0.720512), (13895,-0.781769), (13896,-0.571293), (13897,-0.736136), (13898,-0.764876), (13899,-0.513061), (13900,-0.532051), (13901,-0.686205), (13902,-0.750718), (13903,-0.919268), (13904,-0.656307), (13905,-0.806749), (13906,-0.809940), (13907,-0.565564), (13908,-0.420580), (13909,-0.602605), (13910,-0.627168), (13911,-0.704686), (13912,-0.524868), (13913,-0.719898), (13914,-0.783014), (13915,-0.527486), (13916,-0.522319), (13917,-0.673223), (13918,-0.682451), (13919,-0.854258), (13920,-0.590834), (13921,-0.772859), (13922,-0.811354), (13923,-0.593916), (13924,-0.402488), (13925,-0.550607), (13926,-0.618826), (13927,-0.668010), (13928,-0.577840), (13929,-0.748250), (13930,-0.425371), (13931,-0.569770), (13932,-0.563676), (13933,-0.753133), (13934,-0.869204), (13935,-0.984806), (13936,-0.711163), (13937,-0.906657), (13938,-0.562870), (13939,-0.705416), (13940,-0.576693), (13941,-0.747109), (13942,-0.720570), (13943,-0.873335), (13944,-0.528622), (13945,-0.675813), (13946,-0.722204), (13947,-0.468536), (13948,-0.482410), (13949,-0.614273), (13950,-0.649982), (13951,-0.850585), (13952,-0.754843), (13953,-0.884846), (13954,-0.965144), (13955,-0.726804), (13956,-0.583216), (13957,-0.699750), (13958,-0.771689), (13959,-0.836195), (13960,-0.971771), (13961,-0.687446), (13962,-0.851819), (13963,-0.483418), (13964,-0.672876), (13965,-0.647270), (13966,-0.828369), (13967,-0.870114), (13968,-1.036347), (13969,-0.775710), (13970,-0.942406), (13971,-0.624631), (13972,-0.736519), (13973,-0.580395), (13974,-0.739196), (13975,-0.722413), (13976,-1.000592), (13977,-0.732985), (13978,-0.860202), (13979,-0.548933), (13980,-0.711446), (13981,-0.671445), (13982,-0.840002), (13983,-0.917050), (13984,-1.049839), (13985,-0.825432), (13986,-0.974014), (13987,-0.644629), (13988,-0.789955), (13989,-0.601314), (13990,-0.756865), (13991,-0.747521), (13992,-1.130207), (13993,-0.850985), (13994,-0.611249), (13995,-0.666932), (13996,-0.819233), (13997,-0.810816), (13998,-0.991445), (13999,-1.030873), (14000,-1.192923), (14001,-0.919744), (14002,-0.721811), (14003,-0.751483), (14004,-0.907027), (14005,-0.759263), (14006,-0.827488), (14007,-0.869703), (14008,-1.091671), (14009,-0.815705), (14010,-0.980542), (14011,-0.606568), (14012,-0.770942), (14013,-0.756025), (14014,-0.932007), (14015,-1.004416), (14016,-1.166930), (14017,-0.906755), (14018,-1.059983), (14019,-0.713880), (14020,-0.884290), (14021,-0.724446), (14022,-0.883710), (14023,-0.849745), (14024,-1.018765), (14025,-0.742799), (14026,-0.881162), (14027,-0.537845), (14028,-0.693859), (14029,-0.697984), (14030,-0.853065), (14031,-0.906425), (14032,-1.097743), (14033,-0.803192), (14034,-0.970358), (14035,-0.587556), (14036,-0.768184), (14037,-0.662692), (14038,-0.773184), (14039,-0.738756), (14040,-1.037830), (14041,-0.796704), (14042,-0.934597), (14043,-0.596853), (14044,-0.706882), (14045,-0.706830), (14046,-0.890245), (14047,-0.964507), (14048,-1.146532), (14049,-0.836196), (14050,-0.978272), (14051,-0.630772), (14052,-0.809084), (14053,-0.658063), (14054,-0.811291), (14055,-0.799624), (14056,-0.929627), (14057,-0.668057), (14058,-0.797127), (14059,-0.469602), (14060,-0.610751), (14061,-0.604657), (14062,-0.738373), (14063,-0.820068), (14064,-0.962150), (14065,-0.685250), (14066,-0.840801), (14067,-0.509563), (14068,-0.675327), (14069,-0.476004), (14070,-0.675681), (14071,-0.606412), (14072,-0.904097), (14073,-0.647172), (14074,-0.759524), (14075,-0.443615), (14076,-0.624707), (14077,-0.617686), (14078,-0.779273), (14079,-0.879082), (14080,-1.010476), (14081,-0.721967), (14082,-0.890524), (14083,-0.544421), (14084,-0.691606), (14085,-0.515970), (14086,-0.698459), (14087,-0.675646), (14088,-0.964038), (14089,-0.699218), (14090,-0.860342), (14091,-0.507733), (14092,-0.672106), (14093,-0.651147), (14094,-0.814130), (14095,-0.862381), (14096,-0.997494), (14097,-0.732210), (14098,-0.860817), (14099,-0.523536), (14100,-0.667008), (14101,-0.532713), (14102,-0.726817), (14103,-0.711430), (14104,-0.539044), (14105,-0.696918), (14106,-0.733554), (14107,-0.870526), (14108,-0.442671), (14109,-0.574991), (14110,-0.665977), (14111,-0.797371), (14112,-0.569250), (14113,-0.741056), (14114,-0.790234), (14115,-0.908158), (14116,-0.394837), (14117,-0.529017), (14118,-0.599565), (14119,-0.763006), (14120,-0.596663), (14121,-0.744318), (14122,-0.745186), (14123,-0.495695), (14124,-0.488674), (14125,-0.651651), (14126,-0.705481), (14127,-0.913517), (14128,-0.628259), (14129,-0.796351), (14130,-0.853888), (14131,-0.605330), (14132,-0.442700), (14133,-0.607073), (14134,-0.656251), (14135,-0.714257), (14136,-0.627337), (14137,-0.763377), (14138,-0.810237), (14139,-0.536594), (14140,-0.558365), (14141,-0.728781), (14142,-0.804439), (14143,-0.981354), (14144,-0.692376), (14145,-0.846068), (14146,-0.896178), (14147,-0.647150), (14148,-0.491952), (14149,-0.660509), (14150,-0.719905), (14151,-0.793240), (14152,-0.624111), (14153,-0.768973), (14154,-0.824657), (14155,-0.605359), (14156,-0.564424), (14157,-0.745986), (14158,-0.810029), (14159,-0.994840), (14160,-0.729093), (14161,-0.867919), (14162,-0.951010), (14163,-0.702445), (14164,-0.534706), (14165,-0.683287), (14166,-0.762195), (14167,-0.796514), (14168,-0.479208), (14169,-0.626393), (14170,-0.682540), (14171,-0.816726), (14172,-0.406053), (14173,-0.555567), (14174,-0.605671), (14175,-0.770045), (14176,-0.489902), (14177,-0.636161), (14178,-0.715532), (14179,-0.900807), (14180,-0.339177), (14181,-0.485436), (14182,-0.523931), (14183,-0.673909), (14184,-0.635761), (14185,-0.823822), (14186,-0.475859), (14187,-0.632807), (14188,-0.636462), (14189,-0.777147), (14190,-0.837940), (14191,-0.987449), (14192,-0.718915), (14193,-0.878642), (14194,-0.551118), (14195,-0.731290), (14196,-0.563080), (14197,-0.697730), (14198,-0.667948), (14199,-0.829998), (14200,-0.629742), (14201,-0.746276), (14202,-0.809856), (14203,-0.569187), (14204,-0.526399), (14205,-0.692169), (14206,-0.769217), (14207,-0.964711), (14208,-0.811374), (14209,-0.956236), (14210,-0.993804), (14211,-0.741526), (14212,-0.604444), (14213,-0.748842), (14214,-0.783161), (14215,-0.853240), (14216,-0.979067), (14217,-0.702167), (14218,-0.815915), (14219,-0.504183), (14220,-0.661587), (14221,-0.647597), (14222,-0.798501), (14223,-0.858825), (14224,-1.019948), (14225,-0.786718), (14226,-0.927404), (14227,-0.602196), (14228,-0.765179), (14229,-0.590934), (14230,-0.763210), (14231,-0.723202), (14232,-1.067799), (14233,-0.783937), (14234,-0.944597), (14235,-0.639371), (14236,-0.777733), (14237,-0.769316), (14238,-0.910928), (14239,-0.981940), (14240,-1.096145), (14241,-0.841544), (14242,-0.980376), (14243,-0.679789), (14244,-0.837663), (14245,-0.674100), (14246,-0.846839), (14247,-0.798936), (14248,-0.972601), (14249,-0.687343), (14250,-0.880520), (14251,-0.536271), (14252,-0.685316), (14253,-0.668539), (14254,-0.849631), (14255,-0.924826), (14256,-1.050646), (14257,-0.747736), (14258,-0.936267), (14259,-0.616638), (14260,-0.755928), (14261,-0.629064), (14262,-0.780896), (14263,-0.712097), (14264,-1.069236), (14265,-0.773759), (14266,-0.924663), (14267,-0.587383), (14268,-0.742934), (14269,-0.731730), (14270,-0.886348), (14271,-0.947141), (14272,-1.123593), (14273,-0.843908), (14274,-0.972984), (14275,-0.637094), (14276,-0.781962), (14277,-0.639307), (14278,-0.761408), (14279,-0.769252), (14280,-0.942912), (14281,-0.659513), (14282,-0.862909), (14283,-0.514477), (14284,-0.644943), (14285,-0.622131), (14286,-0.753987), (14287,-0.870058), (14288,-1.052547), (14289,-0.761252), (14290,-0.904261), (14291,-0.575803), (14292,-0.710916), (14293,-0.522275), (14294,-0.680142), (14295,-0.669402), (14296,-1.112013), (14297,-0.846729), (14298,-0.988805), (14299,-0.622264), (14300,-0.768986), (14301,-0.774501), (14302,-0.916119), (14303,-0.994557), (14304,-1.142212), (14305,-0.863923), (14306,-1.011578), (14307,-0.669651), (14308,-0.829842), (14309,-0.696016), (14310,-0.845061), (14311,-0.822242), (14312,-0.965250), (14313,-0.658627), (14314,-0.791880), (14315,-0.476898), (14316,-0.618510), (14317,-0.617988), (14318,-0.780972), (14319,-0.877525), (14320,-1.026576), (14321,-0.765469), (14322,-0.911264), (14323,-0.537754), (14324,-0.716993), (14325,-0.591056), (14326,-0.736851), (14327,-0.728897), (14328,-0.766002), (14329,-0.497469), (14330,-0.639545), (14331,-0.705910), (14332,-0.444346), (14333,-0.422460), (14334,-0.614235), (14335,-0.731696), (14336,-1.123211), (14337,-1.305237), (14338,-1.012545), (14339,-0.767700), (14340,-0.826633), (14341,-0.945954), (14342,-0.791220), (14343,-0.854799), (14344,-1.097206), (14345,-1.284340), (14346,-1.005125), (14347,-0.743554), (14348,-0.764404), (14349,-0.913449), (14350,-0.913391), (14351,-1.076838), (14352,-1.150173), (14353,-1.326155), (14354,-1.054835), (14355,-0.803020), (14356,-0.844772), (14357,-1.016578), (14358,-0.881819), (14359,-0.931923), (14360,-1.062389), (14361,-0.772028), (14362,-0.917353), (14363,-0.972110), (14364,-0.749092), (14365,-0.728603), (14366,-0.845594), (14367,-0.949123), (14368,-1.158086), (14369,-0.895588), (14370,-1.039524), (14371,-1.100317), (14372,-0.845722), (14373,-0.714213), (14374,-0.872543), (14375,-0.941232), (14376,-1.175286), (14377,-0.902570), (14378,-1.037213), (14379,-0.696219), (14380,-0.822966), (14381,-0.792721), (14382,-0.945015), (14383,-1.035539), (14384,-1.181797), (14385,-0.936488), (14386,-1.072991), (14387,-0.725492), (14388,-0.902407), (14389,-0.731881), (14390,-0.899974), (14391,-0.876228), (14392,-1.232435), (14393,-0.975517), (14394,-1.106446), (14395,-0.751978), (14396,-0.934003), (14397,-0.950206), (14398,-1.075094), (14399,-1.160508), (14400,-1.292828), (14401,-1.010825), (14402,-1.132933), (14403,-0.811907), (14404,-0.980927), (14405,-0.806218), (14406,-0.930185), (14407,-0.873459), (14408,-1.150242), (14409,-0.898891), (14410,-1.036790), (14411,-0.723667), (14412,-0.855524), (14413,-0.879154), (14414,-1.003584), (14415,-1.090851), (14416,-1.219458), (14417,-0.952784), (14418,-1.115298), (14419,-0.802639), (14420,-0.925673), (14421,-0.805315), (14422,-0.964579), (14423,-0.908780), (14424,-1.015558), (14425,-0.725654), (14426,-0.925331), (14427,-1.009811), (14428,-0.796556), (14429,-0.745403), (14430,-0.898631), (14431,-0.932943), (14432,-1.104749), (14433,-0.825070), (14434,-1.012204), (14435,-1.051626), (14436,-0.812823), (14437,-0.674808), (14438,-0.828036), (14439,-0.894401), (14440,-1.284984), (14441,-0.978361), (14442,-0.729802), (14443,-0.787802), (14444,-0.955895), (14445,-0.936796), (14446,-1.124394), (14447,-1.179144), (14448,-1.346774), (14449,-1.065698), (14450,-0.823639), (14451,-0.876999), (14452,-1.065061), (14453,-0.935411), (14454,-1.007813), (14455,-1.045845), (14456,-1.271533), (14457,-0.981171), (14458,-1.104668), (14459,-0.749273), (14460,-0.904354), (14461,-0.876432), (14462,-1.046841), (14463,-1.102061), (14464,-1.432726), (14465,-1.147931), (14466,-0.887757), (14467,-0.959702), (14468,-1.110137), (14469,-0.958659), (14470,-1.023628), (14471,-1.076062), (14472,-1.215351), (14473,-1.337459), (14474,-0.720087), (14475,-0.893753), (14476,-0.933638), (14477,-1.078043), (14478,-1.076126), (14479,-1.228427), (14480,-1.306865), (14481,-1.442904), (14482,-0.763292), (14483,-0.937891), (14484,-0.985672), (14485,-1.124968), (14486,-0.907060), (14487,-1.092335), (14488,-1.384910), (14489,-1.534424), (14490,-0.865031), (14491,-1.001070), (14492,-1.075332), (14493,-1.243888), (14494,-1.225715), (14495,-1.378473), (14496,-1.442523), (14497,-1.577166), (14498,-0.850177), (14499,-1.000149), (14500,-1.040041), (14501,-1.183976), (14502,-0.970714), (14503,-1.133234), (14504,-1.226074), (14505,-1.400667), (14506,-0.705263), (14507,-0.878465), (14508,-0.915564), (14509,-1.073901), (14510,-1.062234), (14511,-1.220102), (14512,-1.264176), (14513,-1.450841), (14514,-0.749401), (14515,-0.908201), (14516,-0.967598), (14517,-1.136154), (14518,-0.876443), (14519,-1.034781), (14520,-1.260932), (14521,-1.404404), (14522,-0.739193), (14523,-0.912853), (14524,-0.972719), (14525,-1.147312), (14526,-1.163515), (14527,-1.280043), (14528,-1.361274), (14529,-1.516825), (14530,-0.842322), (14531,-0.970929), (14532,-1.027539), (14533,-1.164975), (14534,-0.933135), (14535,-1.107727), (14536,-1.201964), (14537,-1.373307), (14538,-0.658391), (14539,-0.833447), (14540,-0.895167), (14541,-1.044212), (14542,-1.046946), (14543,-1.188559), (14544,-1.264217), (14545,-1.429980), (14546,-0.751764), (14547,-0.885481), (14548,-0.923513), (14549,-1.090672), (14550,-0.898782), (14551,-1.004627), (14552,-1.305098), (14553,-1.462046), (14554,-0.770355), (14555,-0.931942), (14556,-0.998771), (14557,-1.147816), (14558,-1.137539), (14559,-1.328856), (14560,-1.352956), (14561,-1.502001), (14562,-0.868374), (14563,-1.027638), (14564,-1.077279), (14565,-1.218898), (14566,-0.998203), (14567,-1.138425), (14568,-1.169488), (14569,-1.364982), (14570,-0.719277), (14571,-0.866005), (14572,-0.947229), (14573,-1.084665), (14574,-1.111551), (14575,-1.293576), (14576,-1.337644), (14577,-1.469038), (14578,-0.805687), (14579,-0.983993), (14580,-1.007165), (14581,-1.120907), (14582,-0.864916), (14583,-1.011638), (14584,-0.988818), (14585,-1.161557), (14586,-0.870263), (14587,-0.629594), (14588,-0.690850), (14589,-0.832932), (14590,-0.801753), (14591,-0.980992), (14592,-1.065936), (14593,-1.214518), (14594,-0.943198), (14595,-0.711358), (14596,-0.762858), (14597,-0.893325), (14598,-0.727909), (14599,-0.815639), (14600,-1.001384), (14601,-1.157862), (14602,-0.875853), (14603,-0.650982), (14604,-0.715488), (14605,-0.860820), (14606,-0.838934), (14607,-1.016313), (14608,-1.094288), (14609,-1.276782), (14610,-0.984091), (14611,-0.711375), (14612,-0.773564), (14613,-0.949547), (14614,-0.806429), (14615,-0.856069), (14616,-1.094299), (14617,-0.841094), (14618,-1.020333), (14619,-0.685376), (14620,-0.826525), (14621,-0.822754), (14622,-0.981091), (14623,-1.076718), (14624,-1.217866), (14625,-0.946547), (14626,-1.078403), (14627,-0.743909), (14628,-0.867876), (14629,-0.717789), (14630,-0.897954), (14631,-0.871422), (14632,-1.265717), (14633,-0.969783), (14634,-0.727254), (14635,-0.783870), (14636,-0.945458), (14637,-0.935180), (14638,-1.144143), (14639,-1.173816), (14640,-1.338653), (14641,-1.043645), (14642,-0.818774), (14643,-0.856342), (14644,-1.030002), (14645,-0.875268), (14646,-0.957432), (14647,-1.035407), (14648,-1.135680), (14649,-0.883402), (14650,-1.035239), (14651,-0.716537), (14652,-0.858149), (14653,-0.790278), (14654,-0.982058), (14655,-1.073972), (14656,-1.209548), (14657,-0.942405), (14658,-1.103528), (14659,-0.752779), (14660,-0.900897), (14661,-0.747553), (14662,-0.911927), (14663,-0.880748), (14664,-1.089254), (14665,-0.807709), (14666,-0.981375), (14667,-0.634339), (14668,-0.780134), (14669,-0.768930), (14670,-0.917975), (14671,-1.019181), (14672,-1.194237), (14673,-0.923380), (14674,-1.044554), (14675,-0.677086), (14676,-0.813126), (14677,-0.680690), (14678,-0.886866), (14679,-0.856151), (14680,-1.135720), (14681,-0.823988), (14682,-0.991617), (14683,-0.658050), (14684,-0.797809), (14685,-0.776386), (14686,-0.921248), (14687,-0.999693), (14688,-1.171499), (14689,-0.880204), (14690,-1.035285), (14691,-0.673854), (14692,-0.831728), (14693,-0.708114), (14694,-0.858086), (14695,-0.831090), (14696,-1.063284), (14697,-1.226261), (14698,-0.518778), (14699,-0.667823), (14700,-0.760669), (14701,-0.936652), (14702,-0.948209), (14703,-1.060561), (14704,-1.125067), (14705,-1.278758), (14706,-0.634913), (14707,-0.771415), (14708,-0.831745), (14709,-1.006337), (14710,-0.773571), (14711,-0.908683), (14712,-1.256530), (14713,-0.980101), (14714,-0.714354), (14715,-0.771890), (14716,-0.922795), (14717,-0.936676), (14718,-1.088507), (14719,-1.142331), (14720,-1.525950), (14721,-1.257880), (14722,-1.020467), (14723,-1.040384), (14724,-1.194069), (14725,-1.032372), (14726,-1.091305), (14727,-1.183219), (14728,-1.337373), (14729,-1.025640), (14730,-0.777545), (14731,-0.847161), (14732,-1.001315), (14733,-0.993831), (14734,-1.175856), (14735,-1.222247), (14736,-1.405662), (14737,-1.123196), (14738,-0.861626), (14739,-0.927992), (14740,-1.079360), (14741,-0.894902), (14742,-0.980773), (14743,-1.036456), (14744,-1.289551), (14745,-1.424201), (14746,-0.769666), (14747,-0.925680), (14748,-0.961852), (14749,-1.131805), (14750,-1.143826), (14751,-1.334674), (14752,-1.374565), (14753,-1.515251), (14754,-0.850034), (14755,-1.021840), (14756,-1.074274), (14757,-1.191271), (14758,-0.972900), (14759,-1.135414), (14760,-1.271923), (14761,-1.393561), (14762,-0.717198), (14763,-0.868566), (14764,-0.922859), (14765,-1.110921), (14766,-1.087638), (14767,-1.249225), (14768,-1.329066), (14769,-1.474392), (14770,-0.804072), (14771,-0.941501), (14772,-1.017159), (14773,-1.156918), (14774,-0.929724), (14775,-1.082482), (14776,-1.389923), (14777,-1.533858), (14778,-0.871434), (14779,-1.013510), (14780,-1.080339), (14781,-1.230780), (14782,-1.254880), (14783,-1.398815), (14784,-1.436847), (14785,-1.575209), (14786,-0.909066), (14787,-1.075299), (14788,-1.117977), (14789,-1.301862), (14790,-1.106252), (14791,-1.262729), (14792,-1.258489), (14793,-1.401497), (14794,-0.735354), (14795,-0.899264), (14796,-0.958667), (14797,-1.085414), (14798,-1.110904), (14799,-1.301288), (14800,-1.338856), (14801,-1.489298), (14802,-0.779028), (14803,-0.950834), (14804,-0.984683), (14805,-1.113760), (14806,-0.876347), (14807,-1.066268), (14808,-1.379744), (14809,-1.510674), (14810,-0.838495), (14811,-0.978717), (14812,-1.037650), (14813,-1.176939), (14814,-1.187570), (14815,-1.362163), (14816,-1.434565), (14817,-1.552026), (14818,-0.852439), (14819,-1.026104), (14820,-1.089684), (14821,-1.276355), (14822,-1.045442), (14823,-1.171725), (14824,-1.245987), (14825,-1.384350), (14826,-0.720066), (14827,-0.861215), (14828,-0.915045), (14829,-1.058517), (14830,-1.071928), (14831,-1.192175), (14832,-1.261328), (14833,-1.399227), (14834,-0.708469), (14835,-0.867269), (14836,-0.912264), (14837,-1.086857), (14838,-0.874991), (14839,-0.997562), (14840,-0.966847), (14841,-1.178602), (14842,-0.909136), (14843,-0.623884), (14844,-0.662842), (14845,-0.849977), (14846,-0.816938), (14847,-1.005006), (14848,-1.063476), (14849,-1.230636), (14850,-0.944914), (14851,-0.731189), (14852,-0.777580), (14853,-0.954496), (14854,-0.805804), (14855,-0.855445), (14856,-1.048623), (14857,-1.200917), (14858,-0.921238), (14859,-0.695898), (14860,-0.726960), (14861,-0.881121), (14862,-0.891745), (14863,-1.057045), (14864,-1.113662), (14865,-1.292901), (14866,-1.005782), (14867,-0.753968), (14868,-0.811511), (14869,-0.936868), (14870,-0.768202), (14871,-0.874974), (14872,-1.161976), (14873,-0.885547), (14874,-1.045274), (14875,-0.688025), (14876,-0.837997), (14877,-0.854200), (14878,-1.012068), (14879,-1.084007), (14880,-1.217729), (14881,-0.959878), (14882,-1.115886), (14883,-0.779539), (14884,-0.929047), (14885,-0.745052), (14886,-0.903853), (14887,-0.891253), (14888,-1.298560), (14889,-1.004010), (14890,-0.736409), (14891,-0.809738), (14892,-0.945777), (14893,-0.984742), (14894,-1.162121), (14895,-1.211768), (14896,-1.351058), (14897,-1.078341), (14898,-0.846038), (14899,-0.871527), (14900,-1.052626), (14901,-0.910897), (14902,-0.979123), (14903,-1.009722), (14904,-1.116964), (14905,-0.813591), (14906,-0.971458), (14907,-0.693639), (14908,-0.823172), (14909,-0.824047), (14910,-0.963800), (14911,-1.043171), (14912,-1.208478), (14913,-0.962236), (14914,-1.111750), (14915,-0.787939), (14916,-0.931411), (14917,-0.791079), (14918,-0.915039), (14919,-0.877825), (14920,-1.138346), (14921,-0.880032), (14922,-1.062520), (14923,-0.680187), (14924,-0.814830), (14925,-0.820815), (14926,-1.017705), (14927,-1.105899), (14928,-1.285601), (14929,-0.975265), (14930,-1.108981), (14931,-0.797248), (14932,-0.929575), (14933,-0.782273), (14934,-0.922959), (14935,-0.877842), (14936,-1.168564), (14937,-0.886555), (14938,-1.000766), (14939,-0.664876), (14940,-0.808348), (14941,-0.771596), (14942,-0.916002), (14943,-1.011165), (14944,-1.150454), (14945,-0.869842), (14946,-1.036538), (14947,-0.695081), (14948,-0.866424), (14949,-0.731665), (14950,-0.863522), (14951,-0.829093), (14952,-1.197378), (14953,-0.938600), (14954,-0.725339), (14955,-0.808429), (14956,-0.972340), (14957,-0.973672), (14958,-1.094852), (14959,-1.154249), (14960,-1.326055), (14961,-1.043583), (14962,-0.778769), (14963,-0.824233), (14964,-0.981174), (14965,-0.846878), (14966,-0.883514), (14967,-0.947556), (14968,-1.342785), (14969,-1.071929), (14970,-0.812688), (14971,-0.888803), (14972,-1.028098), (14973,-1.043832), (14974,-1.214712), (14975,-1.254603), (14976,-1.370668), (14977,-1.490915), (14978,-0.830345), (14979,-0.995651), (14980,-1.037396), (14981,-1.197593), (14982,-0.957857), (14983,-1.106902), (14984,-1.262453), (14985,-1.411498), (14986,-0.722130), (14987,-0.880467), (14988,-0.945900), (14989,-1.080549), (14990,-1.112545), (14991,-1.254620), (14992,-1.336315), (14993,-1.477927), (14994,-0.825722), (14995,-0.998455), (14996,-1.044382), (14997,-1.175782), (14998,-0.973666), (14999,-1.103206), (15000,-1.269903), (15001,-1.321866), (15002,-1.093283), (15003,-0.767148), (15004,-0.931058), (15005,-1.000210), (15006,-1.156688), (15007,-1.154776), (15008,-1.295925), (15009,-1.373437), (15010,-1.117446), (15011,-0.829401), (15012,-0.947788), (15013,-1.022983), (15014,-1.100031), (15015,-0.966199), (15016,-1.373970), (15017,-1.098467), (15018,-1.233117), (15019,-0.969686), (15020,-1.110835), (15021,-1.210181), (15022,-1.388957), (15023,-1.352669), (15024,-1.518439), (15025,-1.181158), (15026,-1.309302), (15027,-1.056097), (15028,-1.171235), (15029,-1.138196), (15030,-1.277955), (15031,-1.169207), (15032,-1.330325), (15033,-1.364180), (15034,-1.105396), (15035,-0.807601), (15036,-0.976621), (15037,-1.026262), (15038,-1.224079), (15039,-1.178505), (15040,-1.333123), (15041,-1.386020), (15042,-1.177404), (15043,-0.872641), (15044,-1.041660), (15045,-1.081082), (15046,-1.163710), (15047,-0.997824), (15048,-1.199824), (15049,-1.267586), (15050,-1.051538), (15051,-0.777431), (15052,-0.920903), (15053,-0.957539), (15054,-1.145137), (15055,-1.125110), (15056,-1.274618), (15057,-1.323796), (15058,-1.086846), (15059,-0.787656), (15060,-0.978973), (15061,-1.057418), (15062,-1.125637), (15063,-0.952325), (15064,-1.252332), (15065,-1.270853), (15066,-1.037623), (15067,-0.743078), (15068,-0.959474), (15069,-1.010047), (15070,-1.172561), (15071,-1.134883), (15072,-1.327591), (15073,-1.392560), (15074,-1.151434), (15075,-0.828555), (15076,-0.993856), (15077,-1.075550), (15078,-1.148885), (15079,-1.003437), (15080,-1.152489), (15081,-1.198416), (15082,-0.966576), (15083,-0.661813), (15084,-0.840582), (15085,-0.876290), (15086,-1.039737), (15087,-1.050362), (15088,-1.236106), (15089,-1.291326), (15090,-1.017214), (15091,-0.737998), (15092,-0.919559), (15093,-0.980352), (15094,-1.038822), (15095,-0.879442), (15096,-1.165511), (15097,-1.193787), (15098,-0.972636), (15099,-0.722681), (15100,-0.926997), (15101,-0.975248), (15102,-1.153560), (15103,-1.138174), (15104,-1.258885), (15105,-1.303422), (15106,-1.061363), (15107,-0.745911), (15108,-0.920040), (15109,-0.976187), (15110,-1.030480), (15111,-0.875746), (15112,-1.254714), (15113,-1.308544), (15114,-1.020035), (15115,-0.756605), (15116,-0.900547), (15117,-0.974808), (15118,-1.150791), (15119,-1.155379), (15120,-1.329045), (15121,-1.335493), (15122,-1.140810), (15123,-0.830473), (15124,-0.987877), (15125,-1.053780), (15126,-1.131761), (15127,-0.933365), (15128,-1.210611), (15129,-1.350364), (15130,-0.692586), (15131,-0.814687), (15132,-0.870370), (15133,-1.051469), (15134,-1.042588), (15135,-1.178627), (15136,-1.250566), (15137,-1.416336), (15138,-0.759478), (15139,-0.902487), (15140,-0.960030), (15141,-1.111862), (15142,-0.862840), (15143,-1.018384), (15144,-1.086146), (15145,-1.245410), (15146,-0.559762), (15147,-0.712983), (15148,-0.767276), (15149,-0.959984), (15150,-0.981754), (15151,-1.123836), (15152,-1.161868), (15153,-1.328564), (15154,-0.645239), (15155,-0.793351), (15156,-0.868546), (15157,-1.005975), (15158,-0.751844), (15159,-0.907858), (15160,-1.169312), (15161,-1.349014), (15162,-0.676835), (15163,-0.818910), (15164,-0.888526), (15165,-1.016206), (15166,-1.052378), (15167,-1.226977), (15168,-1.296593), (15169,-1.390829), (15170,-0.728399), (15171,-0.873267), (15172,-0.947992), (15173,-1.108653), (15174,-0.876349), (15175,-1.028644), (15176,-1.188371), (15177,-1.352751), (15178,-0.684748), (15179,-0.829616), (15180,-0.894122), (15181,-1.004614), (15182,-0.999447), (15183,-1.163820), (15184,-1.228332), (15185,-1.385737), (15186,-0.710307), (15187,-0.862602), (15188,-0.909463), (15189,-1.084982), (15190,-0.860574), (15191,-1.025411), (15192,-1.141482), (15193,-1.299350), (15194,-0.681985), (15195,-0.836139), (15196,-0.892286), (15197,-1.033435), (15198,-1.050565), (15199,-1.214476), (15200,-1.286878), (15201,-1.404339), (15202,-0.721007), (15203,-0.848224), (15204,-0.941533), (15205,-1.091968), (15206,-0.841550), (15207,-1.012893), (15208,-1.316613), (15209,-1.039721), (15210,-0.761431), (15211,-0.923945), (15212,-0.968483), (15213,-1.122637), (15214,-1.106324), (15215,-1.246546), (15216,-1.311052), (15217,-1.051805), (15218,-0.788844), (15219,-0.947182), (15220,-0.976391), (15221,-1.065981), (15222,-0.919606), (15223,-1.080730), (15224,-1.155919), (15225,-1.310073), (15226,-0.633254), (15227,-0.788798), (15228,-0.863060), (15229,-1.010715), (15230,-1.023199), (15231,-1.163421), (15232,-1.450423), (15233,-1.511210), (15234,-1.249646), (15235,-0.974143), (15236,-1.158491), (15237,-1.204882), (15238,-1.311661), (15239,-1.142995), (15240,-1.365890), (15241,-1.449907), (15242,-1.225500), (15243,-0.941174), (15244,-1.100902), (15245,-1.143116), (15246,-1.335824), (15247,-1.296286), (15248,-1.479701), (15249,-1.508447), (15250,-1.289612), (15251,-0.970447), (15252,-1.124601), (15253,-1.160773), (15254,-1.246187), (15255,-1.113281), (15256,-1.224706), (15257,-1.294785), (15258,-1.452196), (15259,-0.779553), (15260,-0.905373), (15261,-0.981025), (15262,-1.140289), (15263,-1.157889), (15264,-1.339444), (15265,-1.381196), (15266,-1.545569), (15267,-0.851092), (15268,-0.985741), (15269,-1.046997), (15270,-1.184896), (15271,-0.952123), (15272,-1.270709), (15273,-1.338471), (15274,-1.123350), (15275,-0.861322), (15276,-0.999685), (15277,-1.052582), (15278,-1.242503), (15279,-1.260560), (15280,-1.403569), (15281,-1.466678), (15282,-1.258533), (15283,-0.952373), (15284,-1.123715), (15285,-1.145022), (15286,-1.225790), (15287,-1.071983), (15288,-1.504838), (15289,-1.538224), (15290,-1.300347), (15291,-1.020662), (15292,-1.195254), (15293,-1.236542), (15294,-1.428786), (15295,-1.379493), (15296,-1.522495), (15297,-1.567496), (15298,-1.351918), (15299,-1.057830), (15300,-1.201772), (15301,-1.240730), (15302,-1.332180), (15303,-1.211817), (15304,-1.398952), (15305,-1.439770), (15306,-1.177272), (15307,-0.903166), (15308,-1.081008), (15309,-1.109754), (15310,-1.315931), (15311,-1.322378), (15312,-1.446339), (15313,-1.494590), (15314,-1.266933), (15315,-0.996539), (15316,-1.175315), (15317,-1.190122), (15318,-1.247659), (15319,-1.096181), (15320,-1.264731), (15321,-1.326920), (15322,-1.501976), (15323,-0.812608), (15324,-0.933319), (15325,-0.993649), (15326,-1.177070), (15327,-1.199773), (15328,-1.353928), (15329,-1.420294), (15330,-1.549364), (15331,-0.860929), (15332,-1.038308), (15333,-1.081912), (15334,-1.251395), (15335,-1.039993), (15336,-1.055264), (15337,-1.186664), (15338,-1.244200), (15339,-1.017470), (15340,-0.731754), (15341,-0.872903), (15342,-0.920684), (15343,-1.098996), (15344,-1.090116), (15345,-1.281897), (15346,-1.326891), (15347,-1.089478), (15348,-0.798647), (15349,-0.953271), (15350,-1.003375), (15351,-1.092502), (15352,-1.084085), (15353,-1.120727), (15354,-1.296246), (15355,-0.592019), (15356,-0.749423), (15357,-0.794888), (15358,-0.958798), (15359,-0.991257), (15360,-1.115217), (15361,-1.195515), (15362,-1.357572), (15363,-0.681673), (15364,-0.853942), (15365,-0.920308), (15366,-1.087474), (15367,-0.816611), (15368,-1.033013), (15369,-1.215502), (15370,-1.263289), (15371,-1.047704), (15372,-0.754550), (15373,-0.920783), (15374,-0.988545), (15375,-1.147809), (15376,-1.117094), (15377,-1.296796), (15378,-1.300458), (15379,-1.071867), (15380,-0.800548), (15381,-0.948666), (15382,-1.006203), (15383,-1.070715), (15384,-1.229979), (15385,-1.424083), (15386,-1.136965), (15387,-0.856816), (15388,-0.893457), (15389,-1.085702), (15390,-1.066602), (15391,-1.232365), (15392,-1.292695), (15393,-1.458928), (15394,-1.169024), (15395,-0.910246), (15396,-0.940845), (15397,-1.092676), (15398,-0.933303), (15399,-1.021960), (15400,-1.112483), (15401,-1.167697), (15402,-1.320925), (15403,-0.658501), (15404,-0.798253), (15405,-0.893886), (15406,-1.003451), (15407,-1.036837), (15408,-1.197491), (15409,-1.257821), (15410,-1.421267), (15411,-0.734222), (15412,-0.897206), (15413,-0.965425), (15414,-1.124226), (15415,-0.863588), (15416,-1.107391), (15417,-1.246217), (15418,-0.962355), (15419,-0.752349), (15420,-0.802923), (15421,-0.979369), (15422,-0.966775), (15423,-1.111637), (15424,-1.165461), (15425,-1.364211), (15426,-1.071057), (15427,-0.812742), (15428,-0.854024), (15429,-1.026293), (15430,-0.880852), (15431,-0.952327), (15432,-1.113914), (15433,-1.184000), (15434,-1.327472), (15435,-0.632994), (15436,-0.776003), (15437,-0.864197), (15438,-0.997913), (15439,-1.019226), (15440,-1.176167), (15441,-1.272727), (15442,-1.435704), (15443,-0.769097), (15444,-0.888881), (15445,-0.959430), (15446,-1.084787), (15447,-0.871525), (15448,-1.210549), (15449,-1.358204), (15450,-1.066446), (15451,-0.823454), (15452,-0.880997), (15453,-1.022609), (15454,-1.001650), (15455,-1.136299), (15456,-1.191519), (15457,-1.374934), (15458,-1.086889), (15459,-0.860159), (15460,-0.896337), (15461,-1.066747), (15462,-0.894825), (15463,-0.977452), (15464,-1.165050), (15465,-1.226307), (15466,-0.987497), (15467,-0.690630), (15468,-0.886593), (15469,-0.902791), (15470,-1.136374), (15471,-1.113092), (15472,-1.277465), (15473,-1.336405), (15474,-1.096669), (15475,-0.808160), (15476,-0.956742), (15477,-0.994774), (15478,-1.041165), (15479,-0.892004), (15480,-1.342041), (15481,-1.427455), (15482,-1.197468), (15483,-0.879236), (15484,-1.052438), (15485,-1.102543), (15486,-1.269703), (15487,-1.265468), (15488,-1.620747), (15489,-1.687583), (15490,-1.412544), (15491,-1.125895), (15492,-1.299091), (15493,-1.312039), (15494,-1.400239), (15495,-1.234823), (15496,-1.498131), (15497,-1.559857), (15498,-1.320584), (15499,-1.042295), (15500,-1.185303), (15501,-1.217762), (15502,-1.416043), (15503,-1.407162), (15504,-1.570602), (15505,-1.597025), (15506,-1.355429), (15507,-1.066458), (15508,-1.247086), (15509,-1.329251), (15510,-1.436956), (15511,-1.255741), (15512,-1.363916), (15513,-1.410771), (15514,-1.558889), (15515,-0.871844), (15516,-1.016713), (15517,-1.061707), (15518,-1.239086), (15519,-1.264112), (15520,-1.390403), (15521,-1.431684), (15522,-1.588162), (15523,-0.932237), (15524,-1.084075), (15525,-1.143935), (15526,-1.305522), (15527,-1.071359), (15528,-1.392731), (15529,-1.442842), (15530,-1.189637), (15531,-0.940608), (15532,-1.122633), (15533,-1.186213), (15534,-1.342227), (15535,-1.307799), (15536,-1.486104), (15537,-1.560372), (15538,-1.292766), (15539,-1.031658), (15540,-1.168168), (15541,-1.200157), (15542,-1.294857), (15543,-1.107149), (15544,-1.518170), (15545,-1.583602), (15546,-1.380566), (15547,-1.086948), (15548,-1.222055), (15549,-1.287494), (15550,-1.469519), (15551,-1.414189), (15552,-1.601787), (15553,-1.683482), (15554,-1.412625), (15555,-1.133403), (15556,-1.283844), (15557,-1.341387), (15558,-1.416112), (15559,-1.269275), (15560,-1.438294), (15561,-1.510696), (15562,-1.280716), (15563,-0.972703), (15564,-1.154264), (15565,-1.189040), (15566,-1.350627), (15567,-1.353362), (15568,-1.521912), (15569,-1.571096), (15570,-1.322531), (15571,-1.016840), (15572,-1.172848), (15573,-1.246647), (15574,-1.300940), (15575,-1.149919), (15576,-1.373747), (15577,-1.418748), (15578,-1.607743), (15579,-0.935563), (15580,-1.051628), (15581,-1.120780), (15582,-1.267502), (15583,-1.280919), (15584,-1.462017), (15585,-1.502836), (15586,-1.659313), (15587,-1.000602), (15588,-1.144538), (15589,-1.175600), (15590,-1.335797), (15591,-1.139724), (15592,-1.163817), (15593,-1.343056), (15594,-1.391770), (15595,-1.158540), (15596,-0.884897), (15597,-1.056239), (15598,-1.072437), (15599,-1.257248), (15600,-1.225606), (15601,-1.413668), (15602,-1.462388), (15603,-1.236584), (15604,-0.939253), (15605,-1.105017), (15606,-1.137476), (15607,-1.221493), (15608,-1.269744), (15609,-1.317995), (15610,-1.462857), (15611,-0.784178), (15612,-0.900242), (15613,-0.986583), (15614,-1.132841), (15615,-1.119778), (15616,-1.184754), (15617,-1.255759), (15618,-1.407597), (15619,-0.722875), (15620,-0.903967), (15621,-0.991704), (15622,-1.146785), (15623,-0.913555), (15624,-1.083965), (15625,-1.291074), (15626,-1.347221), (15627,-1.077755), (15628,-0.817117), (15629,-0.939224), (15630,-1.010700), (15631,-1.190865), (15632,-1.199173), (15633,-1.304555), (15634,-1.368134), (15635,-1.177171), (15636,-0.900741), (15637,-1.080907), (15638,-1.128694), (15639,-1.196450), (15640,-1.346428), (15641,-1.529843), (15642,-1.239012), (15643,-1.002068), (15644,-1.015943), (15645,-1.193322), (15646,-1.172832), (15647,-1.355784), (15648,-1.369664), (15649,-1.533568), (15650,-1.244596), (15651,-1.009506), (15652,-1.072159), (15653,-1.219344), (15654,-1.040459), (15655,-1.118904), (15656,-1.207098), (15657,-1.259531), (15658,-1.413686), (15659,-0.749402), (15660,-0.900770), (15661,-0.952734), (15662,-1.130113), (15663,-1.147243), (15664,-1.301867), (15665,-1.331070), (15666,-1.477792), (15667,-0.814905), (15668,-0.982528), (15669,-1.016847), (15670,-1.150100), (15671,-0.921046), (15672,-1.158813), (15673,-1.335728), (15674,-1.063475), (15675,-0.828385), (15676,-0.851552), (15677,-1.017785), (15678,-0.988003), (15679,-1.163522), (15680,-1.243357), (15681,-1.396121), (15682,-1.129911), (15683,-0.899924), (15684,-0.942602), (15685,-1.108835), (15686,-0.934596), (15687,-1.009785), (15688,-1.185310), (15689,-1.227519), (15690,-1.351016), (15691,-0.678373), (15692,-0.831137), (15693,-0.906326), (15694,-1.055834), (15695,-1.076220), (15696,-1.249417), (15697,-1.308813), (15698,-1.449499), (15699,-0.783825), (15700,-0.921724), (15701,-0.988090), (15702,-1.122733), (15703,-0.863492), (15704,-1.215985), (15705,-1.352951), (15706,-1.053297), (15707,-0.832609), (15708,-0.899438), (15709,-1.099578), (15710,-1.065613), (15711,-1.219304), (15712,-1.273128), (15713,-1.434252), (15714,-1.152706), (15715,-0.927372), (15716,-0.999774), (15717,-1.183659), (15718,-1.020566), (15719,-1.088328), (15720,-1.242019), (15721,-1.292123), (15722,-1.036132), (15723,-0.782464), (15724,-0.927326), (15725,-0.984869), (15726,-1.174790), (15727,-1.173336), (15728,-1.376262), (15729,-1.434269), (15730,-1.162949), (15731,-0.901848), (15732,-1.028595), (15733,-1.072200), (15734,-1.172479), (15735,-1.010312), (15736,-1.415291), (15737,-1.462151), (15738,-1.193618), (15739,-0.904177), (15740,-1.081092), (15741,-1.144208), (15742,-1.307192), (15743,-1.290409), (15744,-1.438527), (15745,-1.507216), (15746,-1.643255), (15747,-0.939492), (15748,-1.103865), (15749,-1.168835), (15750,-1.314167), (15751,-1.075357), (15752,-1.327062), (15753,-1.406897), (15754,-1.530394), (15755,-0.882366), (15756,-1.042099), (15757,-1.085704), (15758,-1.247291), (15759,-1.259775), (15760,-1.417179), (15761,-1.486332), (15762,-1.606579), (15763,-0.941832), (15764,-1.103419), (15765,-1.170248), (15766,-1.321616), (15767,-1.072131), (15768,-1.432983), (15769,-1.486807), (15770,-1.620993), (15771,-0.967855), (15772,-1.101108), (15773,-1.176296), (15774,-1.341603), (15775,-1.356873), (15776,-1.483627), (15777,-1.560675), (15778,-1.713433), (15779,-1.045900), (15780,-1.175903), (15781,-1.232976), (15782,-1.386204), (15783,-1.158083), (15784,-1.314561), (15785,-1.353519), (15786,-1.504424), (15787,-0.835031), (15788,-0.984076), (15789,-1.053228), (15790,-1.206456), (15791,-1.215227), (15792,-1.381454), (15793,-1.414376), (15794,-1.605230), (15795,-0.926081), (15796,-1.070016), (15797,-1.122913), (15798,-1.276604), (15799,-1.041515), (15800,-1.374496), (15801,-1.418570), (15802,-1.583407), (15803,-0.925629), (15804,-1.073741), (15805,-1.128035), (15806,-1.284975), (15807,-1.314178), (15808,-1.465553), (15809,-1.528662), (15810,-1.667958), (15811,-0.991595), (15812,-1.152256), (15813,-1.221871), (15814,-1.395537), (15815,-1.120034), (15816,-1.287194), (15817,-1.303392), (15818,-1.498429), (15819,-0.796982), (15820,-0.936741), (15821,-1.025861), (15822,-1.166084), (15823,-1.184610), (15824,-1.357806), (15825,-1.390729), (15826,-1.523055), (15827,-0.855985), (15828,-1.020358), (15829,-1.058853), (15830,-1.206508), (15831,-0.999746), (15832,-1.407517), (15833,-1.463200), (15834,-1.619215), (15835,-0.957717), (15836,-1.127200), (15837,-1.158263), (15838,-1.299882), (15839,-1.320262), (15840,-1.451655), (15841,-1.490613), (15842,-1.647097), (15843,-1.047378), (15844,-1.219184), (15845,-1.289263), (15846,-1.416016), (15847,-1.146549), (15848,-1.201770), (15849,-1.358710), (15850,-1.410674), (15851,-1.138891), (15852,-0.900082), (15853,-1.054706), (15854,-1.107133), (15855,-1.283585), (15856,-1.279814), (15857,-1.409817), (15858,-1.445989), (15859,-1.204394), (15860,-0.920532), (15861,-1.071436), (15862,-1.132229), (15863,-1.195809), (15864,-1.205506), (15865,-1.251434), (15866,-1.398619), (15867,-0.755700), (15868,-0.903818), (15869,-0.950209), (15870,-1.079286), (15871,-1.109422), (15872,-1.262649), (15873,-1.332265), (15874,-1.460872), (15875,-0.778010), (15876,-0.939134), (15877,-1.032437), (15878,-1.177305), (15879,-0.943606), (15880,-1.135850), (15881,-1.334594), (15882,-1.362876), (15883,-1.112921), (15884,-0.824413), (15885,-0.981817), (15886,-1.021245), (15887,-1.204197), (15888,-1.197639), (15889,-1.331356), (15890,-1.408867), (15891,-1.172851), (15892,-0.894561), (15893,-1.068691), (15894,-1.093717), (15895,-1.176801), (15896,-1.092674), (15897,-1.236146), (15898,-0.958320), (15899,-1.107829), (15900,-0.764512), (15901,-0.923313), (15902,-0.914895), (15903,-1.076482), (15904,-1.140988), (15905,-1.270528), (15906,-0.993629), (15907,-1.140357), (15908,-0.796571), (15909,-0.969773), (15910,-0.813180), (15911,-0.978950), (15912,-1.226466), (15913,-1.248242), (15914,-1.450705), (15915,-0.764124), (15916,-0.932680), (15917,-0.997186), (15918,-1.156914), (15919,-1.163825), (15920,-1.283146), (15921,-1.346262), (15922,-1.482764), (15923,-0.858893), (15924,-1.004219), (15925,-1.066408), (15926,-1.191765), (15927,-0.930658), (15928,-1.207441), (15929,-1.369961), (15930,-1.110250), (15931,-0.842644), (15932,-0.894614), (15933,-1.094284), (15934,-1.061252), (15935,-1.259996), (15936,-1.268767), (15937,-1.428031), (15938,-1.170180), (15939,-0.904896), (15940,-0.987054), (15941,-1.142605), (15942,-0.993907), (15943,-1.062596), (15944,-1.229293), (15945,-1.285440), (15946,-1.462355), (15947,-0.790639), (15948,-0.932721), (15949,-0.981898), (15950,-1.121194), (15951,-1.122063), (15952,-1.272504), (15953,-1.332827), (15954,-1.475373), (15955,-0.815272), (15956,-0.971286), (15957,-1.018604), (15958,-1.186233), (15959,-0.967862), (15960,-1.036087), (15961,-1.225076), (15962,-0.956542), (15963,-1.109770), (15964,-0.769703), (15965,-0.941046), (15966,-0.922873), (15967,-1.083533), (15968,-1.139680), (15969,-1.272000), (15970,-1.009039), (15971,-1.167376), (15972,-0.781324), (15973,-0.943844), (15974,-0.811865), (15975,-0.994823), (15976,-1.170342), (15977,-1.218130), (15978,-1.360675), (15979,-0.701501), (15980,-0.826858), (15981,-0.906229), (15982,-1.071066), (15983,-1.075654), (15984,-1.224236), (15985,-1.279919), (15986,-1.467517), (15987,-0.775826), (15988,-0.920695), (15989,-0.987060), (15990,-1.143538), (15991,-0.903339), (15992,-1.222388), (15993,-1.266926), (15994,-1.398782), (15995,-0.724279), (15996,-0.889116), (15997,-0.928081), (15998,-1.094778), (15999,-1.100756), (16000,-1.508527), (16001,-1.547955), (16002,-1.275239), (16003,-1.035503), (16004,-1.172005), (16005,-1.229549), (16006,-1.319139), (16007,-1.154186), (16008,-1.318096), (16009,-1.469464), (16010,-1.114069), (16011,-1.286801), (16012,-1.014085), (16013,-1.192861), (16014,-1.245294), (16015,-1.406418), (16016,-1.395208), (16017,-1.522425), (16018,-1.203722), (16019,-1.367633), (16020,-1.088880), (16021,-1.255577), (16022,-1.223008), (16023,-1.370193), (16024,-1.203850), (16025,-1.338493), (16026,-1.393250), (16027,-1.153051), (16028,-0.864542), (16029,-1.018697), (16030,-1.132902), (16031,-1.316787), (16032,-1.283755), (16033,-1.422581), (16034,-1.478727), (16035,-1.222266), (16036,-0.922149), (16037,-1.110674), (16038,-1.141743), (16039,-1.238296), (16040,-1.288406), (16041,-1.436525), (16042,-1.066727), (16043,-1.232497), (16044,-0.933307), (16045,-1.104186), (16046,-1.206782), (16047,-1.340498), (16048,-1.338580), (16049,-1.504814), (16050,-1.142455), (16051,-1.282208), (16052,-1.017388), (16053,-1.172012), (16054,-1.184032), (16055,-1.317749), (16056,-1.419881), (16057,-1.546628), (16058,-1.231182), (16059,-1.396483), (16060,-1.104725), (16061,-1.247733), (16062,-1.331751), (16063,-1.506807), (16064,-1.522077), (16065,-1.653940), (16066,-1.330129), (16067,-1.444340), (16068,-1.159545), (16069,-1.302553), (16070,-1.284380), (16071,-1.471052), (16072,-1.372986), (16073,-1.556401), (16074,-1.192646), (16075,-1.317540), (16076,-1.031818), (16077,-1.211057), (16078,-1.277886), (16079,-1.426004), (16080,-1.401795), (16081,-1.551767), (16082,-1.194981), (16083,-1.348672), (16084,-1.073170), (16085,-1.239403), (16086,-1.205901), (16087,-1.345191), (16088,-1.234589), (16089,-1.405462), (16090,-1.454176), (16091,-1.209331), (16092,-0.926402), (16093,-1.074983), (16094,-1.138563), (16095,-1.308972), (16096,-1.334462), (16097,-1.491872), (16098,-1.556842), (16099,-1.309210), (16100,-1.034170), (16101,-1.179502), (16102,-1.237972), (16103,-1.308521), (16104,-1.136599), (16105,-1.268455), (16106,-1.351083), (16107,-1.078366), (16108,-0.770347), (16109,-0.937513), (16110,-0.993196), (16111,-1.196123), (16112,-1.192345), (16113,-1.345573), (16114,-1.384068), (16115,-1.143405), (16116,-0.871153), (16117,-1.052251), (16118,-1.089356), (16119,-1.151076), (16120,-1.037681), (16121,-1.181617), (16122,-1.241946), (16123,-0.958084), (16124,-0.722525), (16125,-0.897117), (16126,-0.919820), (16127,-1.116711), (16128,-1.163102), (16129,-1.299611), (16130,-1.352971), (16131,-1.120668), (16132,-0.819154), (16133,-0.994210), (16134,-1.011804), (16135,-1.118119), (16136,-1.112951), (16137,-1.270819), (16138,-1.309784), (16139,-1.029635), (16140,-0.755992), (16141,-0.912469), (16142,-0.985804), (16143,-1.167360), (16144,-1.140364), (16145,-1.303348), (16146,-1.345093), (16147,-1.103497), (16148,-0.833110), (16149,-0.982155), (16150,-1.022973), (16151,-1.104204), (16152,-1.266718), (16153,-1.335870), (16154,-1.473306), (16155,-0.787188), (16156,-0.962713), (16157,-1.030469), (16158,-1.159076), (16159,-1.172956), (16160,-1.297850), (16161,-1.362356), (16162,-1.525803), (16163,-0.866629), (16164,-1.003595), (16165,-1.059742), (16166,-1.222725), (16167,-1.015969), (16168,-1.221219), (16169,-1.275506), (16170,-1.444989), (16171,-0.761200), (16172,-0.907922), (16173,-0.979861), (16174,-1.122406), (16175,-1.138603), (16176,-1.302977), (16177,-1.380025), (16178,-1.507242), (16179,-0.830416), (16180,-0.948340), (16181,-0.994268), (16182,-1.173043), (16183,-0.927734), (16184,-1.178037), (16185,-1.215142), (16186,-1.368833), (16187,-0.700366), (16188,-0.832693), (16189,-0.888839), (16190,-1.034171), (16191,-1.059661), (16192,-1.223571), (16193,-1.276005), (16194,-1.424580), (16195,-0.753797), (16196,-0.912134), (16197,-0.957598), (16198,-1.099210), (16199,-0.896631), (16200,-1.139044), (16201,-1.209586), (16202,-1.354918), (16203,-0.665550), (16204,-0.820637), (16205,-0.893040), (16206,-1.049054), (16207,-1.053642), (16208,-1.220802), (16209,-1.230499), (16210,-1.404629), (16211,-0.735699), (16212,-0.888927), (16213,-0.950646), (16214,-1.113166), (16215,-0.865534), (16216,-1.210131), (16217,-1.266278), (16218,-1.434834), (16219,-0.762655), (16220,-0.914023), (16221,-0.972023), (16222,-1.101563), (16223,-1.095468), (16224,-1.261232), (16225,-1.315062), (16226,-1.452491), (16227,-0.765446), (16228,-0.927503), (16229,-1.040781), (16230,-1.193076), (16231,-0.964956), (16232,-1.238019), (16233,-1.265832), (16234,-1.028419), (16235,-0.751989), (16236,-0.927978), (16237,-0.964150), (16238,-1.118768), (16239,-1.110814), (16240,-1.288663), (16241,-1.359205), (16242,-1.135261), (16243,-0.841180), (16244,-0.983262), (16245,-1.034762), (16246,-1.140608), (16247,-0.981234), (16248,-1.381566), (16249,-1.428427), (16250,-1.165003), (16251,-0.910402), (16252,-1.055734), (16253,-1.140678), (16254,-1.344531), (16255,-1.299420), (16256,-1.055038), (16257,-1.188755), (16258,-0.846371), (16259,-0.979624), (16260,-0.713877), (16261,-0.867562), (16262,-0.819201), (16263,-1.000300), (16264,-0.963079), (16265,-1.115843), (16266,-0.783209), (16267,-0.958265), (16268,-0.696700), (16269,-0.840636), (16270,-0.919544), (16271,-1.044901), (16272,-1.037873), (16273,-1.201784), (16274,-0.862643), (16275,-0.983361), (16276,-0.704138), (16277,-0.855043), (16278,-0.820151), (16279,-0.958977), (16280,-0.885532), (16281,-1.068021), (16282,-0.715412), (16283,-0.851915), (16284,-0.579668), (16285,-0.774229), (16286,-0.868002), (16287,-1.000329), (16288,-1.003984), (16289,-1.144206), (16290,-0.810645), (16291,-0.968049), (16292,-0.685114), (16293,-0.820227), (16294,-0.819705), (16295,-0.962251), (16296,-1.039299), (16297,-0.825574), (16298,-0.891476), (16299,-1.034485), (16300,-0.741794), (16301,-0.926142), (16302,-0.972070), (16303,-1.123438), (16304,-1.115020), (16305,-0.878071), (16306,-0.955582), (16307,-1.153869), (16308,-0.890445), (16309,-0.963774), (16310,-1.011098), (16311,-1.144814), (16312,-1.031420), (16313,-1.212519), (16314,-0.843191), (16315,-1.014064), (16316,-0.738098), (16317,-0.877857), (16318,-0.970234), (16319,-1.086298), (16320,-1.082527), (16321,-1.236682), (16322,-0.906834), (16323,-1.021972), (16324,-0.744609), (16325,-0.897837), (16326,-0.846220), (16327,-0.998521), (16328,-0.873981), (16329,-1.043464), (16330,-0.694569), (16331,-0.842687), (16332,-0.582976), (16333,-0.750606), (16334,-0.832763), (16335,-0.986918), (16336,-0.980823), (16337,-1.124296), (16338,-0.795374), (16339,-0.949066), (16340,-0.675423), (16341,-0.821681), (16342,-0.779820), (16343,-0.927938), (16344,-0.966433), (16345,-1.134990), (16346,-0.798636), (16347,-0.961156), (16348,-0.682397), (16349,-0.821229), (16350,-0.896418), (16351,-1.041286), (16352,-1.057484), (16353,-1.220467), (16354,-0.863212), (16355,-0.974167), (16356,-0.718639), (16357,-0.872793), (16358,-0.854157), (16359,-1.022713), (16360,-0.855901), (16361,-0.909731), (16362,-0.673244), (16363,-0.751689), (16364,-0.900271), (16365,-0.603866), (16366,-0.782172), (16367,-0.826710), (16368,-0.991083), (16369,-0.997062), (16370,-0.763368), (16371,-0.812545), (16372,-0.940689), (16373,-0.640102), (16374,-0.708791), (16375,-0.759365), (16376,-0.870326), (16377,-1.020761), (16378,-0.666762), (16379,-0.795369), (16380,-0.546341), (16381,-0.687959), (16382,-0.768721), (16383,-0.924271), (16384,-0.907031), (16385,-1.066295), (16386,-0.739697), (16387,-0.904071), (16388,-0.636001), (16389,-0.733024), (16390,-0.705565), (16391,-0.862505), (16392,-0.856875), (16393,-0.919058), (16394,-0.707192), (16395,-0.762876), (16396,-0.918890), (16397,-0.623876), (16398,-0.786859), (16399,-0.834647), (16400,-0.990191), (16401,-0.979451), (16402,-0.739715), (16403,-0.803764), (16404,-0.963028), (16405,-0.674056), (16406,-0.749244), (16407,-0.810964), (16408,-0.985093), (16409,-1.035204), (16410,-0.793145), (16411,-0.530647), (16412,-0.681089), (16413,-0.722834), (16414,-0.898823), (16415,-0.909910), (16416,-1.058492), (16417,-1.092347), (16418,-0.865617), (16419,-0.587791), (16420,-0.774925), (16421,-0.831535), (16422,-0.920199), (16423,-0.748740), (16424,-0.832294), (16425,-1.004564), (16426,-0.654278), (16427,-0.782891), (16428,-0.497169), (16429,-0.593259), (16430,-0.677740), (16431,-0.856052), (16432,-0.838342), (16433,-0.996680), (16434,-0.648717), (16435,-0.801945), (16436,-0.537588), (16437,-0.687566), (16438,-0.671716), (16439,-0.828657), (16440,-1.008822), (16441,-1.046854), (16442,-0.816873), (16443,-0.500494), (16444,-0.662081), (16445,-0.708942), (16446,-0.909082), (16447,-0.893232), (16448,-1.080830), (16449,-1.129545), (16450,-0.861938), (16451,-0.592014), (16452,-0.733163), (16453,-0.785127), (16454,-0.876577), (16455,-0.710698), (16456,-0.860206), (16457,-1.026439), (16458,-0.693805), (16459,-0.826595), (16460,-0.566884), (16461,-0.726148), (16462,-0.781368), (16463,-0.944345), (16464,-0.916886), (16465,-1.074753), (16466,-0.721218), (16467,-0.872122), (16468,-0.629137), (16469,-0.787004), (16470,-0.759545), (16471,-0.906267), (16472,-0.981462), (16473,-1.015774), (16474,-0.766282), (16475,-0.472664), (16476,-0.630538), (16477,-0.681576), (16478,-0.864997), (16479,-0.840318), (16480,-0.978217), (16481,-1.028791), (16482,-0.791842), (16483,-0.517272), (16484,-0.695578), (16485,-0.755907), (16486,-0.851534), (16487,-0.659643), (16488,-0.901123), (16489,-0.664173), (16490,-0.703595), (16491,-0.886553), (16492,-0.639848), (16493,-0.834879), (16494,-0.866874), (16495,-0.991298), (16496,-0.996819), (16497,-0.769162), (16498,-0.792792), (16499,-0.953916), (16500,-0.675626), (16501,-0.760571), (16502,-0.785133), (16503,-0.978768), (16504,-0.855624), (16505,-0.998626), (16506,-0.672498), (16507,-0.802501), (16508,-0.518633), (16509,-0.685799), (16510,-0.754018), (16511,-0.918398), (16512,-1.026104), (16513,-1.071098), (16514,-0.824863), (16515,-0.700323), (16516,-0.841008), (16517,-0.889722), (16518,-0.979776), (16519,-0.696377), (16520,-1.044694), (16521,-1.059031), (16522,-0.802113), (16523,-0.819243), (16524,-1.004518), (16525,-1.043014), (16526,-1.210173), (16527,-0.908196), (16528,-1.079539), (16529,-1.126394), (16530,-0.933576), (16531,-0.757941), (16532,-0.885151), (16533,-0.903678), (16534,-0.943563), (16535,-0.642049), (16536,-0.871920), (16537,-1.057658), (16538,-0.711555), (16539,-0.848521), (16540,-0.847537), (16541,-1.013307), (16542,-1.075490), (16543,-1.274240), (16544,-0.953678), (16545,-1.087864), (16546,-0.743151), (16547,-0.897305), (16548,-0.760223), (16549,-0.912988), (16550,-0.899924), (16551,-1.071267), (16552,-0.840353), (16553,-1.010300), (16554,-0.643295), (16555,-0.799773), (16556,-0.809471), (16557,-0.957589), (16558,-1.039283), (16559,-1.182755), (16560,-0.921185), (16561,-1.063267), (16562,-0.718554), (16563,-0.860629), (16564,-0.765820), (16565,-0.873062), (16566,-0.840950), (16567,-1.031341), (16568,-0.898435), (16569,-1.037261), (16570,-0.694871), (16571,-0.831844), (16572,-0.843864), (16573,-0.968288), (16574,-1.077390), (16575,-1.243160), (16576,-0.933750), (16577,-1.100910), (16578,-0.743655), (16579,-0.885267), (16580,-0.764447), (16581,-0.922778), (16582,-0.878130), (16583,-1.021139), (16584,-0.805091), (16585,-0.955996), (16586,-0.612216), (16587,-0.775193), (16588,-0.768635), (16589,-0.934868), (16590,-0.992875), (16591,-1.158175), (16592,-0.865021), (16593,-1.030790), (16594,-0.671682), (16595,-0.816081), (16596,-0.672962), (16597,-0.827580), (16598,-0.830772), (16599,-1.010944), (16600,-0.971406), (16601,-1.113945), (16602,-0.744617), (16603,-0.886693), (16604,-0.867130), (16605,-1.018961), (16606,-1.122953), (16607,-1.265492), (16608,-0.965838), (16609,-1.106061), (16610,-0.799901), (16611,-0.927581), (16612,-0.795608), (16613,-0.945116), (16614,-0.924157), (16615,-1.092713), (16616,-0.826966), (16617,-0.961146), (16618,-0.625262), (16619,-0.745509), (16620,-0.725477), (16621,-0.927940), (16622,-1.068625), (16623,-1.202342), (16624,-0.912907), (16625,-1.096328), (16626,-0.755329), (16627,-0.898337), (16628,-0.754286), (16629,-0.887539), (16630,-0.873085), (16631,-1.049537), (16632,-0.807942), (16633,-0.963956), (16634,-0.576507), (16635,-0.758532), (16636,-0.688337), (16637,-0.860607), (16638,-0.943234), (16639,-1.109931), (16640,-0.862762), (16641,-1.017380), (16642,-0.658271), (16643,-0.812426), (16644,-0.655369), (16645,-0.791871), (16646,-0.801569), (16647,-0.955260), (16648,-0.844189), (16649,-0.990917), (16650,-0.646204), (16651,-0.776207), (16652,-0.757101), (16653,-0.913585), (16654,-1.005492), (16655,-1.176835), (16656,-0.891583), (16657,-1.012757), (16658,-0.669440), (16659,-0.820808), (16660,-0.681403), (16661,-0.850886), (16662,-0.800196), (16663,-0.959930), (16664,-0.759210), (16665,-0.802352), (16666,-0.964865), (16667,-0.549552), (16668,-0.738083), (16669,-0.777968), (16670,-0.939092), (16671,-0.686350), (16672,-0.850724), (16673,-0.900834), (16674,-1.045696), (16675,-0.467811), (16676,-0.641014), (16677,-0.689265), (16678,-0.817408), (16679,-0.436465), (16680,-0.893002), (16681,-0.922674), (16682,-0.696407), (16683,-0.684277), (16684,-0.814743), (16685,-0.888078), (16686,-1.059884), (16687,-0.804350), (16688,-0.984985), (16689,-1.019767), (16690,-0.781421), (16691,-0.624364), (16692,-0.783628), (16693,-0.806801), (16694,-0.904751), (16695,-0.603700), (16696,-0.873977), (16697,-0.927807), (16698,-0.685748), (16699,-0.658283), (16700,-0.824053), (16701,-0.878803), (16702,-1.077090), (16703,-0.816916), (16704,-0.964101), (16705,-1.011425), (16706,-0.770762), (16707,-0.616492), (16708,-0.756244), (16709,-0.809141), (16710,-0.871331), (16711,-0.580963), (16712,-0.841021), (16713,-0.878126), (16714,-0.676943), (16715,-0.682921), (16716,-0.810138), (16717,-0.878827), (16718,-1.081290), (16719,-0.815543), (16720,-0.939503), (16721,-0.985895), (16722,-0.714111), (16723,-0.587711), (16724,-0.752548), (16725,-0.789653), (16726,-0.862525), (16727,-0.575870), (16728,-0.654778), (16729,-0.747155), (16730,-0.914321), (16731,-0.544987), (16732,-0.722836), (16733,-0.766441), (16734,-0.886688), (16735,-0.640909), (16736,-0.811326), (16737,-0.831706), (16738,-1.010481), (16739,-0.489721), (16740,-0.674069), (16741,-0.701882), (16742,-0.826312), (16743,-0.434687), (16744,-0.796472), (16745,-0.853546), (16746,-0.609163), (16747,-0.615611), (16748,-0.744688), (16749,-0.804548), (16750,-0.988896), (16751,-0.703174), (16752,-0.848042), (16753,-0.921835), (16754,-0.664917), (16755,-0.507860), (16756,-0.669447), (16757,-0.748355), (16758,-0.831909), (16759,-0.526212), (16760,-0.825287), (16761,-0.878184), (16762,-0.658422), (16763,-0.648609), (16764,-0.776752), (16765,-0.851484), (16766,-1.040472), (16767,-0.751963), (16768,-0.923306), (16769,-1.071424), (16770,-0.709529), (16771,-0.845106), (16772,-0.728455), (16773,-0.881683), (16774,-0.851901), (16775,-0.990727), (16776,-0.796050), (16777,-0.975282), (16778,-0.633362), (16779,-0.778224), (16780,-0.780489), (16781,-0.915138), (16782,-0.985217), (16783,-1.130549), (16784,-0.850400), (16785,-1.011987), (16786,-0.689109), (16787,-0.829794), (16788,-0.703858), (16789,-0.873810), (16790,-0.840309), (16791,-0.994000), (16792,-0.886178), (16793,-1.018968), (16794,-0.696090), (16795,-0.856744), (16796,-0.846936), (16797,-1.015486), (16798,-1.106010), (16799,-1.243445), (16800,-0.968869), (16801,-1.085867), (16802,-0.765305), (16803,-0.895772), (16804,-0.773092), (16805,-0.947221), (16806,-0.881666), (16807,-1.058581), (16808,-1.129130), (16809,-0.849914), (16810,-0.627360), (16811,-0.665861), (16812,-0.811187), (16813,-0.831103), (16814,-1.020561), (16815,-1.088323), (16816,-1.259666), (16817,-0.987877), (16818,-0.782047), (16819,-0.810793), (16820,-0.973770), (16821,-0.811604), (16822,-0.902591), (16823,-0.913215), (16824,-1.221119), (16825,-0.963731), (16826,-0.719818), (16827,-0.753204), (16828,-0.918974), (16829,-0.901264), (16830,-1.106514), (16831,-1.086018), (16832,-1.260610), (16833,-0.968389), (16834,-0.764883), (16835,-0.801988), (16836,-0.972861), (16837,-0.789793), (16838,-0.850586), (16839,-0.892800), (16840,-1.118025), (16841,-0.825334), (16842,-0.554941), (16843,-0.596692), (16844,-0.771284), (16845,-0.762867), (16846,-0.924917), (16847,-0.946224), (16848,-1.097592), (16849,-0.830918), (16850,-0.554026), (16851,-0.606916), (16852,-0.798697), (16853,-0.643037), (16854,-0.733090), (16855,-0.804102), (16856,-1.217910), (16857,-0.960522), (16858,-0.690592), (16859,-0.710978), (16860,-0.903686), (16861,-0.905951), (16862,-1.097732), (16863,-1.151092), (16864,-1.299667), (16865,-1.023701), (16866,-0.792794), (16867,-0.826643), (16868,-0.989163), (16869,-0.847898), (16870,-0.930056), (16871,-0.981556), (16872,-1.131071), (16873,-0.843953), (16874,-0.620478), (16875,-0.671516), (16876,-0.787117), (16877,-0.796351), (16878,-0.973267), (16879,-1.042883), (16880,-1.228158), (16881,-0.940582), (16882,-0.653001), (16883,-0.723080), (16884,-0.907428), (16885,-0.750377), (16886,-0.787939), (16887,-0.870097), (16888,-0.922531), (16889,-0.659107), (16890,-0.809548), (16891,-0.454616), (16892,-0.606447), (16893,-0.603603), (16894,-0.777269), (16895,-0.838988), (16896,-0.987570), (16897,-0.706494), (16898,-0.865295), (16899,-0.546130), (16900,-0.704004), (16901,-0.559952), (16902,-0.707137), (16903,-0.666209), (16904,-0.993618), (16905,-0.728334), (16906,-0.853691), (16907,-0.526630), (16908,-0.689613), (16909,-0.672837), (16910,-0.834887), (16911,-0.903113), (16912,-1.047048), (16913,-0.764113), (16914,-0.899226), (16915,-0.613040), (16916,-0.773694), (16917,-0.605955), (16918,-0.755933), (16919,-0.741943), (16920,-0.659206), (16921,-0.782240), (16922,-0.824448), (16923,-0.612582), (16924,-0.640859), (16925,-0.773185), (16926,-0.811680), (16927,-0.972804), (16928,-0.665717), (16929,-0.848206), (16930,-0.904816), (16931,-0.662293), (16932,-0.480158), (16933,-0.649178), (16934,-0.687673), (16935,-0.773081), (16936,-0.748871), (16937,-0.908599), (16938,-0.529979), (16939,-0.693889), (16940,-0.697550), (16941,-0.836839), (16942,-0.929216), (16943,-1.095913), (16944,-0.816234), (16945,-1.003368), (16946,-0.640540), (16947,-0.800737), (16948,-0.654363), (16949,-0.783433), (16950,-0.732286), (16951,-0.906415), (16952,-0.591426), (16953,-0.743727), (16954,-0.791045), (16955,-0.558278), (16956,-0.573085), (16957,-0.729100), (16958,-0.763882), (16959,-0.973771), (16960,-0.676440), (16961,-0.849173), (16962,-0.907643), (16963,-0.691131), (16964,-0.542903), (16965,-0.681266), (16966,-0.723011), (16967,-0.797279), (16968,-0.613278), (16969,-0.766969), (16970,-0.815220), (16971,-0.580130), (16972,-0.555457), (16973,-0.720294), (16974,-0.778301), (16975,-0.941278), (16976,-0.643483), (16977,-0.813893), (16978,-0.903947), (16979,-0.668857), (16980,-0.476966), (16981,-0.627408), (16982,-0.699346), (16983,-0.748524), (16984,-0.568706), (16985,-0.709391), (16986,-0.793872), (16987,-0.546704), (16988,-0.544792), (16989,-0.701733), (16990,-0.772282), (16991,-0.944088), (16992,-0.658366), (16993,-0.822276), (16994,-0.845906), (16995,-0.628468), (16996,-0.431468), (16997,-0.599091), (16998,-0.648738), (16999,-0.754584), (17000,-0.706687), (17001,-0.852945), (17002,-0.570936), (17003,-0.719981), (17004,-0.716210), (17005,-0.840171), (17006,-0.895391), (17007,-1.056978), (17008,-0.774512), (17009,-0.952355), (17010,-0.623433), (17011,-0.771552), (17012,-0.600563), (17013,-0.751931), (17014,-0.737477), (17015,-0.860041), (17016,-0.736898), (17017,-0.905448), (17018,-0.537047), (17019,-0.674946), (17020,-0.649810), (17021,-0.785386), (17022,-0.863824), (17023,-1.025881), (17024,-0.963582), (17025,-1.124699), (17026,-0.819009), (17027,-0.945293), (17028,-0.822143), (17029,-0.972121), (17030,-0.934443), (17031,-1.101603), (17032,-0.927357), (17033,-1.075475), (17034,-0.733086), (17035,-0.902569), (17036,-0.874176), (17037,-0.993961), (17038,-1.106312), (17039,-1.254430), (17040,-0.991470), (17041,-1.142838), (17042,-0.801844), (17043,-0.950426), (17044,-0.802655), (17045,-0.974931), (17046,-0.959081), (17047,-1.103479), (17048,-1.107141), (17049,-0.844180), (17050,-0.987183), (17051,-0.656872), (17052,-0.795234), (17053,-0.782171), (17054,-0.924716), (17055,-0.986899), (17056,-1.148486), (17057,-0.877629), (17058,-1.022498), (17059,-0.694510), (17060,-0.855627), (17061,-0.680461), (17062,-0.825787), (17063,-0.800188), (17064,-1.127133), (17065,-0.837228), (17066,-0.613754), (17067,-0.663395), (17068,-0.824982), (17069,-0.811918), (17070,-0.996266), (17071,-1.036158), (17072,-1.207964), (17073,-0.938034), (17074,-0.681580), (17075,-0.768383), (17076,-0.937866), (17077,-0.790102), (17078,-0.844389), (17079,-0.906572), (17080,-1.307374), (17081,-0.981245), (17082,-0.767520), (17083,-0.803692), (17084,-0.967602), (17085,-0.915986), (17086,-1.121705), (17087,-1.182028), (17088,-1.343615), (17089,-1.046284), (17090,-0.828377), (17091,-0.876627), (17092,-1.041934), (17093,-0.889060), (17094,-0.987936), (17095,-1.077063), (17096,-1.279990), (17097,-0.998914), (17098,-0.753605), (17099,-0.785601), (17100,-0.964839), (17101,-0.948056), (17102,-1.129155), (17103,-1.181119), (17104,-1.350139), (17105,-0.991030), (17106,-0.745258), (17107,-0.801404), (17108,-0.962522), (17109,-0.784563), (17110,-0.869514), (17111,-0.907546), (17112,-1.103966), (17113,-0.802453), (17114,-0.962650), (17115,-0.676001), (17116,-0.813894), (17117,-0.813373), (17118,-1.000977), (17119,-1.062233), (17120,-1.204309), (17121,-0.919050), (17122,-1.060199), (17123,-0.722456), (17124,-0.882189), (17125,-0.731169), (17126,-0.873251), (17127,-0.836499), (17128,-0.993440), (17129,-0.752308), (17130,-0.910182), (17131,-0.564542), (17132,-0.704294), (17133,-0.672189), (17134,-0.827270), (17135,-0.921977), (17136,-1.075668), (17137,-0.769044), (17138,-0.947813), (17139,-0.615179), (17140,-0.760048), (17141,-0.617856), (17142,-0.770151), (17143,-0.739435), (17144,-0.938649), (17145,-0.659896), (17146,-0.813587), (17147,-0.475380), (17148,-0.642077), (17149,-0.580705), (17150,-0.756694), (17151,-0.843961), (17152,-0.989756), (17153,-0.719363), (17154,-0.850756), (17155,-0.513939), (17156,-0.682032), (17157,-0.551913), (17158,-0.700031), (17159,-0.667462), (17160,-0.980012), (17161,-0.680815), (17162,-0.855877), (17163,-0.516737), (17164,-0.702012), (17165,-0.691272), (17166,-0.866797), (17167,-0.955461), (17168,-1.101719), (17169,-0.787200), (17170,-0.959006), (17171,-0.612897), (17172,-0.750333), (17173,-0.612787), (17174,-0.751150), (17175,-0.730654), (17176,-0.685543), (17177,-0.813686), (17178,-0.876796), (17179,-0.632883), (17180,-0.606351), (17181,-0.786516), (17182,-0.839877), (17183,-1.024688), (17184,-0.752435), (17185,-0.889871), (17186,-0.952054), (17187,-0.720214), (17188,-0.563627), (17189,-0.702453), (17190,-0.791580), (17191,-0.845867), (17192,-0.676737), (17193,-0.829959), (17194,-0.844766), (17195,-0.592488), (17196,-0.591040), (17197,-0.766096), (17198,-0.816669), (17199,-1.009377), (17200,-0.744563), (17201,-0.881066), (17202,-0.941395), (17203,-0.693763), (17204,-0.583155), (17205,-0.745206), (17206,-0.781841), (17207,-0.849603), (17208,-0.666999), (17209,-0.796539), (17210,-0.881946), (17211,-0.672404), (17212,-0.662590), (17213,-0.816281), (17214,-0.879397), (17215,-1.055386), (17216,-0.776164), (17217,-0.940544), (17218,-0.993904), (17219,-0.745339), (17220,-0.589679), (17221,-0.746156), (17222,-0.783261), (17223,-0.829652), (17224,-0.674918), (17225,-0.817457), (17226,-0.815546), (17227,-0.591138), (17228,-0.597117), (17229,-0.750344), (17230,-0.822283), (17231,-0.988516), (17232,-0.699545), (17233,-0.859742), (17234,-0.896377), (17235,-0.652458), (17236,-0.523742), (17237,-0.727595), (17238,-0.759127), (17239,-0.795763), (17240,-0.610835), (17241,-0.778464), (17242,-0.822532), (17243,-0.577687), (17244,-0.589244), (17245,-0.729930), (17246,-0.782827), (17247,-0.928616), (17248,-0.635931), (17249,-0.786372), (17250,-0.845305), (17251,-0.560047), (17252,-0.440153), (17253,-0.605917), (17254,-0.652777), (17255,-0.729826), (17256,-0.677282), (17257,-0.832827), (17258,-0.502052), (17259,-0.621373), (17260,-0.597627), (17261,-0.755495), (17262,-0.855304), (17263,-1.007135), (17264,-0.747431), (17265,-0.901585), (17266,-0.552226), (17267,-0.716600), (17268,-0.586023), (17269,-0.764329), (17270,-0.728974), (17271,-0.880342), (17272,-0.839871), (17273,-1.000068), (17274,-0.625161), (17275,-0.771890), (17276,-0.742101), (17277,-0.901835), (17278,-0.990955), (17279,-1.160445), (17280,-0.837560), (17281,-0.981495), (17282,-1.060867), (17283,-0.830886), (17284,-0.686371), (17285,-0.832167), (17286,-0.877631), (17287,-0.963972), (17288,-0.752570), (17289,-0.900224), (17290,-0.960548), (17291,-0.710593), (17292,-0.687780), (17293,-0.846111), (17294,-0.880893), (17295,-1.074996), (17296,-0.801817), (17297,-0.951325), (17298,-1.024197), (17299,-0.790034), (17300,-0.618111), (17301,-0.767626), (17302,-0.851174), (17303,-0.936124), (17304,-1.082383), (17305,-0.837537), (17306,-0.979613), (17307,-0.643266), (17308,-0.773726), (17309,-0.765308), (17310,-0.968705), (17311,-1.010450), (17312,-1.171573), (17313,-0.883528), (17314,-1.046975), (17315,-0.694366), (17316,-0.802535), (17317,-0.667776), (17318,-0.827509), (17319,-0.762418), (17320,-1.217101), (17321,-0.941605), (17322,-0.715337), (17323,-0.771948), (17324,-0.935858), (17325,-0.931623), (17326,-1.122471), (17327,-1.146571), (17328,-1.346241), (17329,-1.070745), (17330,-0.832399), (17331,-0.906660), (17332,-1.043163), (17333,-0.894935), (17334,-0.951082), (17335,-0.977968), (17336,-1.157670), (17337,-0.891923), (17338,-1.040968), (17339,-0.708797), (17340,-0.869457), (17341,-0.869399), (17342,-1.007762), (17343,-1.089920), (17344,-1.270085), (17345,-0.972291), (17346,-1.111117), (17347,-0.796598), (17348,-0.972117), (17349,-0.855473), (17350,-0.989659), (17351,-0.931999), (17352,-1.137249), (17353,-0.843631), (17354,-1.027053), (17355,-0.681877), (17356,-0.835104), (17357,-0.803462), (17358,-0.941825), (17359,-1.020263), (17360,-1.147943), (17361,-0.885446), (17362,-1.064685), (17363,-0.694894), (17364,-0.837433), (17365,-0.717539), (17366,-0.830817), (17367,-0.840515), (17368,-1.134023), (17369,-0.841332), (17370,-1.000596), (17371,-0.658669), (17372,-0.814220), (17373,-0.828101), (17374,-0.993401), (17375,-1.050011), (17376,-1.190233), (17377,-0.894762), (17378,-1.063312), (17379,-0.737184), (17380,-0.873686), (17381,-0.723599), (17382,-0.867071), (17383,-0.831709), (17384,-1.006302), (17385,-0.746598), (17386,-0.897033), (17387,-0.558362), (17388,-0.715766), (17389,-0.692020), (17390,-0.819237), (17391,-0.902328), (17392,-1.041154), (17393,-0.775870), (17394,-0.913769), (17395,-0.561160), (17396,-0.709279), (17397,-0.566154), (17398,-0.708699), (17399,-0.676588), (17400,-0.994710), (17401,-0.714568), (17402,-0.904489), (17403,-0.525869), (17404,-0.671194), (17405,-0.686001), (17406,-0.801609), (17407,-0.923247), (17408,-1.089943), (17409,-0.802368), (17410,-0.954663), (17411,-0.607627), (17412,-0.758068), (17413,-0.641887), (17414,-0.764458), (17415,-0.757430), (17416,-1.058371), (17417,-0.787515), (17418,-0.934700), (17419,-0.579304), (17420,-0.719063), (17421,-0.739443), (17422,-0.872233), (17423,-0.954391), (17424,-1.098789), (17425,-0.826536), (17426,-1.008562), (17427,-0.658745), (17428,-0.824509), (17429,-0.685573), (17430,-0.816967), (17431,-0.785788), (17432,-0.736031), (17433,-0.892509), (17434,-0.960734), (17435,-0.716815), (17436,-0.681454), (17437,-0.845834), (17438,-0.856922), (17439,-1.025478), (17440,-0.724891), (17441,-0.905989), (17442,-0.975142), (17443,-0.732156), (17444,-0.554197), (17445,-0.712528), (17446,-0.764962), (17447,-0.867094), (17448,-0.620389), (17449,-0.756428), (17450,-0.818618), (17451,-0.600710), (17452,-0.576037), (17453,-0.745057), (17454,-0.797954), (17455,-0.979509), (17456,-0.700757), (17457,-0.852125), (17458,-0.905022), (17459,-0.655067), (17460,-0.491510), (17461,-0.667029), (17462,-0.705994), (17463,-0.790938), (17464,-0.708665), (17465,-0.861892), (17466,-0.898528), (17467,-0.672730), (17468,-0.699610), (17469,-0.854234), (17470,-0.913630), (17471,-1.061285), (17472,-0.779740), (17473,-0.969198), (17474,-1.049502), (17475,-0.813479), (17476,-0.645740), (17477,-0.791535), (17478,-0.870906), (17479,-0.939132), (17480,-0.736553), (17481,-0.908828), (17482,-0.936641), (17483,-0.715483), (17484,-0.711712), (17485,-0.837069), (17486,-0.904825), (17487,-1.069662), (17488,-0.805775), (17489,-0.963179), (17490,-0.976133), (17491,-0.733140), (17492,-0.579340), (17493,-0.733031), (17494,-0.787318), (17495,-0.860189), (17496,-0.670616), (17497,-0.852177), (17498,-0.896245), (17499,-0.665802), (17500,-0.660171), (17501,-0.798997), (17502,-0.853753), (17503,-1.031596), (17504,-0.734728), (17505,-0.917217), (17506,-0.958968), (17507,-0.726658), (17508,-0.589576), (17509,-0.765101), (17510,-0.805920), (17511,-0.902943), (17512,-0.833674), (17513,-0.988762), (17514,-0.628257), (17515,-0.781015), (17516,-0.790713), (17517,-0.957409), (17518,-1.020062), (17519,-1.150065), (17520,-0.863880), (17521,-1.032900), (17522,-0.692833), (17523,-0.842341), (17524,-0.689930), (17525,-0.858950), (17526,-0.844960), (17527,-0.985176), (17528,-0.708746), (17529,-0.862437), (17530,-0.904652), (17531,-0.663056), (17532,-0.648133), (17533,-0.796251), (17534,-0.873299), (17535,-1.055788), (17536,-0.893158), (17537,-1.034776), (17538,-1.068625), (17539,-0.825176), (17540,-0.687624), (17541,-0.818091), (17542,-0.888176), (17543,-0.956402), (17544,-1.108233), (17545,-0.844809), (17546,-1.001750), (17547,-0.648214), (17548,-0.803295), (17549,-0.829248), (17550,-0.934637), (17551,-1.007966), (17552,-1.176522), (17553,-0.881514), (17554,-1.061680), (17555,-0.723473), (17556,-0.866012), (17557,-0.721960), (17558,-0.900736), (17559,-0.850515), (17560,-1.171424), (17561,-0.859692), (17562,-1.018029), (17563,-0.656127), (17564,-0.811215), (17565,-0.805121), (17566,-0.947196), (17567,-1.044219), (17568,-1.177009), (17569,-0.887104), (17570,-1.053338), (17571,-0.723490), (17572,-0.949641), (17573,-0.767506), (17574,-0.954641), (17575,-0.940644), (17576,-1.353525), (17577,-1.066876), (17578,-0.818311), (17579,-0.845661), (17580,-1.030472), (17581,-0.982575), (17582,-1.175746), (17583,-1.235149), (17584,-1.384657), (17585,-1.071528), (17586,-0.834585), (17587,-0.874470), (17588,-1.040240), (17589,-0.837660), (17590,-0.895203), (17591,-0.956923), (17592,-1.118047), (17593,-0.832788), (17594,-1.010174), (17595,-0.682179), (17596,-0.876283), (17597,-0.831172), (17598,-0.984864), (17599,-1.105111), (17600,-1.236041), (17601,-0.993518), (17602,-1.125375), (17603,-0.795064), (17604,-0.963620), (17605,-0.801917), (17606,-0.970473), (17607,-0.903065), (17608,-1.093449), (17609,-0.836988), (17610,-1.025056), (17611,-0.652472), (17612,-0.793621), (17613,-0.771735), (17614,-0.939358), (17615,-1.034991), (17616,-1.172421), (17617,-0.907137), (17618,-1.053865), (17619,-0.745382), (17620,-0.864233), (17621,-0.730871), (17622,-0.871093), (17623,-0.853383), (17624,-1.191481), (17625,-0.898790), (17626,-1.068273), (17627,-0.705445), (17628,-0.845203), (17629,-0.841432), (17630,-0.995123), (17631,-1.065666), (17632,-1.213321), (17633,-0.939208), (17634,-1.086863), (17635,-0.727284), (17636,-0.896774), (17637,-0.742040), (17638,-0.872507), (17639,-0.858047), (17640,-1.023353), (17641,-0.761319), (17642,-0.902932), (17643,-0.543823), (17644,-0.693331), (17645,-0.669585), (17646,-0.841391), (17647,-0.934701), (17648,-1.091642), (17649,-0.819859), (17650,-0.985159), (17651,-0.672030), (17652,-0.784381), (17653,-0.613856), (17654,-0.785198), (17655,-0.756806), (17656,-1.078179), (17657,-0.798500), (17658,-0.948008), (17659,-0.584253), (17660,-0.714256), (17661,-0.721631), (17662,-0.862316), (17663,-0.987210), (17664,-1.116280), (17665,-0.824059), (17666,-0.975427), (17667,-0.657188), (17668,-0.793228), (17669,-0.659865), (17670,-0.836781), (17671,-0.774945), (17672,-1.075879), (17673,-0.773439), (17674,-0.943849), (17675,-0.591703), (17676,-0.763509), (17677,-0.758348), (17678,-0.914362), (17679,-1.012775), (17680,-1.155784), (17681,-0.885854), (17682,-1.038618), (17683,-0.695765), (17684,-0.889863), (17685,-0.750927), (17686,-0.893466), (17687,-0.860897), (17688,-0.682939), (17689,-0.800863), (17690,-0.876052), (17691,-1.022780), (17692,-0.629758), (17693,-0.800168), (17694,-0.827981), (17695,-0.977032), (17696,-0.724290), (17697,-0.876585), (17698,-0.888142), (17699,-1.039510), (17700,-0.507141), (17701,-0.639468), (17702,-0.725802), (17703,-0.894358), (17704,-0.699681), (17705,-0.858018), (17706,-0.900227), (17707,-0.664673), (17708,-0.605624), (17709,-0.763961), (17710,-0.794097), (17711,-0.971013), (17712,-0.706656), (17713,-0.860810), (17714,-0.944828), (17715,-0.686050), (17716,-0.568473), (17717,-0.723560), (17718,-0.798285), (17719,-0.838177), (17720,-0.806072), (17721,-0.948611), (17722,-0.978747), (17723,-0.741797), (17724,-0.715265), (17725,-0.863846), (17726,-0.926962), (17727,-1.111774), (17728,-0.852996), (17729,-0.969987), (17730,-1.049828), (17731,-0.824951), (17732,-0.659072), (17733,-0.818799), (17734,-0.841502), (17735,-0.918557), (17736,-0.723410), (17737,-0.898929), (17738,-0.956936), (17739,-0.705590), (17740,-0.656297), (17741,-0.835536), (17742,-0.907938), (17743,-1.091823), (17744,-0.807960), (17745,-0.937494), (17746,-1.002470), (17747,-0.755764), (17748,-0.592208), (17749,-0.748216), (17750,-0.810868), (17751,-0.890703), (17752,-0.602195), (17753,-0.742417), (17754,-0.816215), (17755,-0.951328), (17756,-0.552734), (17757,-0.717107), (17758,-0.755139), (17759,-0.917189), (17760,-0.686282), (17761,-0.841827), (17762,-0.911449), (17763,-1.035873), (17764,-0.495144), (17765,-0.667414), (17766,-0.711488), (17767,-0.853100), (17768,-1.139176), (17769,-0.869709), (17770,-0.670386), (17771,-0.716777), (17772,-0.856999), (17773,-0.827674), (17774,-1.037107), (17775,-1.063993), (17776,-1.218610), (17777,-0.941254), (17778,-0.720097), (17779,-0.811077), (17780,-0.986139), (17781,-0.822576), (17782,-0.874547), (17783,-0.918151), (17784,-0.772240), (17785,-0.898993), (17786,-0.961176), (17787,-0.718654), (17788,-0.729278), (17789,-0.863001), (17790,-0.947018), (17791,-1.088631), (17792,-1.216311), (17793,-0.943595), (17794,-1.107505), (17795,-0.770224), (17796,-0.896045), (17797,-0.749670), (17798,-0.899185), (17799,-0.868470), (17800,-1.154539), (17801,-0.880896), (17802,-1.037843), (17803,-0.664332), (17804,-0.873759), (17805,-0.878810), (17806,-1.042720), (17807,-1.112342), (17808,-1.266033), (17809,-1.009572), (17810,-1.151185), (17811,-0.800899), (17812,-0.949950), (17813,-0.824477), (17814,-0.905708), (17815,-0.871743), (17816,-1.162458), (17817,-0.872090), (17818,-1.044366), (17819,-0.683861), (17820,-0.822687), (17821,-0.825415), (17822,-0.980966), (17823,-1.060801), (17824,-1.220065), (17825,-0.922270), (17826,-1.062023), (17827,-0.714987), (17828,-0.910487), (17829,-0.766436), (17830,-0.916877), (17831,-0.875010), (17832,-1.185706), (17833,-1.306880), (17834,-0.615189), (17835,-0.781886), (17836,-0.860794), (17837,-1.007979), (17838,-1.013500), (17839,-1.180660), (17840,-1.213582), (17841,-1.384925), (17842,-0.707173), (17843,-0.852498), (17844,-0.925370), (17845,-1.057226), (17846,-0.842111), (17847,-1.010204), (17848,-1.192229), (17849,-0.916727), (17850,-1.046260), (17851,-0.715486), (17852,-0.840843), (17853,-0.833815), (17854,-0.991226), (17855,-1.103577), (17856,-1.259122), (17857,-0.969224), (17858,-1.129878), (17859,-0.806999), (17860,-0.946758), (17861,-0.805956), (17862,-0.947105), (17863,-0.921506), (17864,-1.012486), (17865,-1.183366), (17866,-0.907400), (17867,-0.675096), (17868,-0.688507), (17869,-0.845448), (17870,-0.873724), (17871,-1.044603), (17872,-1.031077), (17873,-1.188017), (17874,-0.924130), (17875,-0.658846), (17876,-0.714530), (17877,-0.891446), (17878,-0.730675), (17879,-0.824906), (17880,-1.135596), (17881,-0.853130), (17882,-1.021217), (17883,-0.679296), (17884,-0.831128), (17885,-0.805985), (17886,-0.957353), (17887,-1.035335), (17888,-1.164875), (17889,-0.910737), (17890,-1.062105), (17891,-0.731793), (17892,-0.864120), (17893,-0.733537), (17894,-0.898374), (17895,-0.873238), (17896,-0.893618), (17897,-1.044059), (17898,-0.766234), (17899,-0.538107), (17900,-0.613301), (17901,-0.790217), (17902,-0.764148), (17903,-0.939204), (17904,-0.997674), (17905,-1.148578), (17906,-0.901410), (17907,-0.647272), (17908,-0.715961), (17909,-0.891950), (17910,-0.736289), (17911,-0.761779), (17912,-1.059927), (17913,-0.793253), (17914,-0.919537), (17915,-0.615236), (17916,-0.720619), (17917,-0.725207), (17918,-0.845454), (17919,-0.950373), (17920,-1.058542), (17921,-0.795581), (17922,-0.967387), (17923,-0.652405), (17924,-0.790767), (17925,-0.652759), (17926,-0.852899), (17927,-0.774801), (17928,-0.984697), (17929,-1.125846), (17930,-0.859636), (17931,-0.606431), (17932,-0.678370), (17933,-0.836707), (17934,-0.835722), (17935,-0.960610), (17936,-0.992605), (17937,-1.193209), (17938,-0.895878), (17939,-0.665428), (17940,-0.707642), (17941,-0.843682), (17942,-0.685235), (17943,-0.735345), (17944,-0.900182), (17945,-0.606101), (17946,-0.792303), (17947,-0.849846), (17948,-0.617079), (17949,-0.593333), (17950,-0.757243), (17951,-0.759972), (17952,-0.951283), (17953,-0.691578), (17954,-0.845269), (17955,-0.894910), (17956,-0.645888), (17957,-0.482789), (17958,-0.673179), (17959,-0.700522), (17960,-0.927607), (17961,-0.657213), (17962,-0.778388), (17963,-0.444827), (17964,-0.600841), (17965,-0.593350), (17966,-0.743791), (17967,-0.837558), (17968,-0.981030), (17969,-0.710643), (17970,-0.870834), (17971,-0.559565), (17972,-0.699787), (17973,-0.572460), (17974,-0.702457), (17975,-0.651774), (17976,-1.008450), (17977,-0.760354), (17978,-0.941910), (17979,-0.572119), (17980,-0.710018), (17981,-0.704850), (17982,-0.881766), (17983,-0.962997), (17984,-1.101823), (17985,-0.815638), (17986,-0.990694), (17987,-0.615323), (17988,-0.766691), (17989,-0.617073), (17990,-0.751716), (17991,-0.735403), (17992,-1.008936), (17993,-0.703703), (17994,-0.849035), (17995,-0.515937), (17996,-0.695639), (17997,-0.668174), (17998,-0.817219), (17999,-0.902633), (18000,-1.073043), (18001,-0.810082), (18002,-0.947981), (18003,-0.626493), (18004,-0.771361), (18005,-0.646821), (18006,-0.775891), (18007,-0.736353), (18008,-0.894221), (18009,-0.582025), (18010,-0.730606), (18011,-0.802082), (18012,-0.560492), (18013,-0.570190), (18014,-0.686255), (18015,-0.749371), (18016,-0.921640), (18017,-0.654497), (18018,-0.807261), (18019,-0.866194), (18020,-0.658042), (18021,-0.495876), (18022,-0.663042), (18023,-0.708970), (18024,-1.151574), (18025,-0.848201), (18026,-0.594533), (18027,-0.647893), (18028,-0.797864), (18029,-0.819178), (18030,-1.016068), (18031,-1.072215), (18032,-1.210577), (18033,-0.928105), (18034,-0.681400), (18035,-0.716645), (18036,-0.849898), (18037,-0.695634), (18038,-0.777322), (18039,-0.836262), (18040,-1.008068), (18041,-0.729309), (18042,-0.887646), (18043,-0.579633), (18044,-0.719849), (18045,-0.718864), (18046,-0.859550), (18047,-0.915233), (18048,-1.249611), (18049,-0.961103), (18050,-1.120367), (18051,-0.758472), (18052,-0.924242), (18053,-0.778794), (18054,-0.932948), (18055,-0.878551), (18056,-1.140000), (18057,-0.841272), (18058,-0.988464), (18059,-0.635855), (18060,-0.789083), (18061,-0.769513), (18062,-0.957581), (18063,-1.026270), (18064,-1.158126), (18065,-0.912354), (18066,-1.049320), (18067,-0.726442), (18068,-0.897784), (18069,-0.727722), (18070,-0.881413), (18071,-0.842802), (18072,-1.088465), (18073,-1.235650), (18074,-0.961543), (18075,-0.703229), (18076,-0.748693), (18077,-0.929322), (18078,-0.908826), (18079,-1.097357), (18080,-1.142821), (18081,-1.288616), (18082,-1.008468), (18083,-0.767335), (18084,-0.838347), (18085,-1.012940), (18086,-0.837304), (18087,-0.904133), (18088,-0.991407), (18089,-1.151134), (18090,-0.862163), (18091,-0.613134), (18092,-0.675787), (18093,-0.807180), (18094,-0.774142), (18095,-0.956637), (18096,-1.040648), (18097,-1.220820), (18098,-0.916983), (18099,-0.684680), (18100,-0.739893), (18101,-0.923778), (18102,-0.772294), (18103,-0.855385), (18104,-1.046233), (18105,-1.212466), (18106,-0.912349), (18107,-0.687008), (18108,-0.754307), (18109,-0.901955), (18110,-0.871247), (18111,-1.047693), (18112,-1.053677), (18113,-1.232916), (18114,-0.992716), (18115,-0.744621), (18116,-0.802621), (18117,-0.999048), (18118,-0.837345), (18119,-0.886529), (18120,-0.997021), (18121,-1.158608), (18122,-0.867313), (18123,-0.641509), (18124,-0.677218), (18125,-0.822550), (18126,-0.848503), (18127,-1.020772), (18128,-1.067633), (18129,-1.229683), (18130,-0.947681), (18131,-0.658240), (18132,-0.705564), (18133,-0.862968), (18134,-0.742147), (18135,-0.787142), (18136,-1.103875), (18137,-1.245487), (18138,-1.002038), (18139,-0.767875), (18140,-0.808229), (18141,-0.986535), (18142,-0.955357), (18143,-1.148064), (18144,-1.226972), (18145,-1.323532), (18146,-1.029914), (18147,-0.813402), (18148,-0.846788), (18149,-0.984224), (18150,-0.842959), (18151,-0.969712), (18152,-0.997988), (18153,-1.143320), (18154,-0.872927), (18155,-0.645733), (18156,-0.696770), (18157,-0.836992), (18158,-0.820673), (18159,-1.000381), (18160,-1.069997), (18161,-1.247376), (18162,-0.939826), (18163,-0.704729), (18164,-0.736725), (18165,-0.865795), (18166,-0.746828), (18167,-0.823413), (18168,-0.910217), (18169,-1.055085), (18170,-0.757285), (18171,-0.518945), (18172,-0.573232), (18173,-0.763153), (18174,-0.716183), (18175,-0.946053), (18176,-1.002200), (18177,-1.140563), (18178,-0.873882), (18179,-0.611855), (18180,-0.660569), (18181,-0.810541), (18182,-0.670209), (18183,-0.754226), (18184,-0.978518), (18185,-1.151257), (18186,-0.853456), (18187,-0.609074), (18188,-0.667080), (18189,-0.831924), (18190,-0.783557), (18191,-0.988343), (18192,-1.056099), (18193,-1.148945), (18194,-0.883662), (18195,-0.659718), (18196,-0.695890), (18197,-0.850044), (18198,-0.710175), (18199,-0.811845), (18200,-0.921873), (18201,-0.643120), (18202,-0.821889), (18203,-0.878969), (18204,-0.614149), (18205,-0.561606), (18206,-0.725516), (18207,-0.786309), (18208,-0.976693), (18209,-0.688648), (18210,-0.852095), (18211,-0.942612), (18212,-0.694053), (18213,-0.527241), (18214,-0.704156), (18215,-0.748231), (18216,-1.090968), (18217,-0.800137), (18218,-0.963120), (18219,-0.605401), (18220,-0.753056), (18221,-0.749749), (18222,-0.889964), (18223,-0.973055), (18224,-1.148574), (18225,-0.879578), (18226,-1.025373), (18227,-0.662545), (18228,-0.810663), (18229,-0.720957), (18230,-0.908091), (18231,-0.859724), (18232,-1.158805), (18233,-0.862864), (18234,-0.997977), (18235,-0.650014), (18236,-0.796273), (18237,-0.778563), (18238,-0.923432), (18239,-1.017668), (18240,-1.134660), (18241,-0.842438), (18242,-1.006812), (18243,-0.653739), (18244,-0.793962), (18245,-0.624362), (18246,-0.788273), (18247,-0.743625), (18248,-1.006470), (18249,-0.753728), (18250,-0.909742), (18251,-0.563639), (18252,-0.716397), (18253,-0.747930), (18254,-0.919272), (18255,-0.956834), (18256,-1.072442), (18257,-0.776965), (18258,-0.948307), (18259,-0.628215), (18260,-0.787010), (18261,-0.632282), (18262,-0.783650), (18263,-0.816103), (18264,-0.911272), (18265,-0.609289), (18266,-0.762516), (18267,-0.797762), (18268,-0.566855), (18269,-0.558901), (18270,-0.703299), (18271,-0.771062), (18272,-0.917783), (18273,-0.652036), (18274,-0.783893), (18275,-0.824248), (18276,-0.624925), (18277,-0.471117), (18278,-0.630388), (18279,-0.680492), (18280,-1.006047), (18281,-0.740300), (18282,-0.905600), (18283,-0.583185), (18284,-0.725731), (18285,-0.697802), (18286,-0.871468), (18287,-0.937833), (18288,-1.083629), (18289,-0.803943), (18290,-0.942775), (18291,-0.633829), (18292,-0.784264), (18293,-0.611885), (18294,-0.774398), (18295,-0.733928), (18296,-1.020930), (18297,-0.760292), (18298,-0.914910), (18299,-0.564630), (18300,-0.753618), (18301,-0.739165), (18302,-0.927690), (18303,-0.989416), (18304,-1.357700), (18305,-1.063619), (18306,-1.211268), (18307,-0.862378), (18308,-1.003991), (18309,-0.849727), (18310,-1.001558), (18311,-0.969916), (18312,-1.154728), (18313,-0.915918), (18314,-1.034776), (18315,-0.677521), (18316,-0.837711), (18317,-0.824184), (18318,-0.982522), (18319,-1.044241), (18320,-1.214657), (18321,-0.921040), (18322,-1.089126), (18323,-0.730018), (18324,-0.917616), (18325,-0.787966), (18326,-0.943047), (18327,-0.922094), (18328,-1.257399), (18329,-0.973073), (18330,-1.141160), (18331,-0.759290), (18332,-0.947352), (18333,-0.937081), (18334,-1.063365), (18335,-1.151095), (18336,-1.321511), (18337,-0.984694), (18338,-1.107265), (18339,-0.781600), (18340,-0.930181), (18341,-0.804708), (18342,-0.962112), (18343,-0.943946), (18344,-1.025170), (18345,-1.202556), (18346,-0.901969), (18347,-0.644118), (18348,-0.677503), (18349,-0.869284), (18350,-0.880372), (18351,-1.010838), (18352,-1.060022), (18353,-1.228109), (18354,-0.932168), (18355,-0.684073), (18356,-0.727677), (18357,-0.902740), (18358,-0.766121), (18359,-0.838523), (18360,-1.174297), (18361,-1.302440), (18362,-1.027401), (18363,-0.770477), (18364,-0.809905), (18365,-0.975675), (18366,-1.006737), (18367,-1.168788), (18368,-1.201246), (18369,-1.387918), (18370,-1.109629), (18371,-0.872679), (18372,-0.924643), (18373,-1.101559), (18374,-0.931966), (18375,-1.001581), (18376,-0.993627), (18377,-1.129203), (18378,-0.841159), (18379,-0.591203), (18380,-0.629235), (18381,-0.819620), (18382,-0.794947), (18383,-0.951425), (18384,-1.020577), (18385,-1.159403), (18386,-0.890869), (18387,-0.659962), (18388,-0.720285), (18389,-0.873050), (18390,-0.661648), (18391,-0.741946), (18392,-1.078653), (18393,-1.240240), (18394,-0.930831), (18395,-0.718495), (18396,-0.766283), (18397,-0.944125), (18398,-0.936171), (18399,-1.120520), (18400,-1.160874), (18401,-1.288091), (18402,-1.023734), (18403,-0.743128), (18404,-0.813670), (18405,-1.037499), (18406,-0.864650), (18407,-0.915687), (18408,-0.958828), (18409,-1.104160), (18410,-0.843522), (18411,-0.598214), (18412,-0.652037), (18413,-0.813624), (18414,-0.794988), (18415,-1.000701), (18416,-1.041056), (18417,-1.196143), (18418,-0.917391), (18419,-0.737573), (18420,-0.801152), (18421,-0.930685), (18422,-0.745294), (18423,-0.809807), (18424,-0.768873), (18425,-0.885407), (18426,-0.644274), (18427,-0.806325), (18428,-0.474154), (18429,-0.620412), (18430,-0.604563), (18431,-0.790307), (18432,-1.234308), (18433,-0.968091), (18434,-1.125502), (18435,-0.781252), (18436,-0.951205), (18437,-0.805294), (18438,-0.963631), (18439,-0.912478), (18440,-1.104259), (18441,-1.269096), (18442,-0.978264), (18443,-0.720883), (18444,-0.776097), (18445,-0.954872), (18446,-0.960387), (18447,-1.128943), (18448,-1.193919), (18449,-1.358756), (18450,-1.065601), (18451,-0.815646), (18452,-0.836959), (18453,-1.020838), (18454,-0.877719), (18455,-0.976133), (18456,-1.345350), (18457,-1.081926), (18458,-1.230971), (18459,-0.885332), (18460,-1.021834), (18461,-1.031995), (18462,-1.155499), (18463,-1.252052), (18464,-1.428505), (18465,-1.171117), (18466,-1.346179), (18467,-1.002856), (18468,-1.123573), (18469,-0.989278), (18470,-1.123457), (18471,-1.096462), (18472,-1.258049), (18473,-0.987655), (18474,-1.145523), (18475,-0.836577), (18476,-1.007919), (18477,-0.971631), (18478,-1.107207), (18479,-1.199584), (18480,-1.326338), (18481,-1.071736), (18482,-1.228214), (18483,-0.865856), (18484,-1.021863), (18485,-0.858307), (18486,-0.985060), (18487,-0.967814), (18488,-1.217190), (18489,-0.950053), (18490,-1.102811), (18491,-0.766927), (18492,-0.920618), (18493,-0.888976), (18494,-1.044990), (18495,-1.143403), (18496,-1.291058), (18497,-1.025311), (18498,-1.168313), (18499,-0.813387), (18500,-0.988443), (18501,-0.840679), (18502,-1.005052), (18503,-0.971551), (18504,-1.215817), (18505,-0.924059), (18506,-1.086573), (18507,-0.761834), (18508,-0.874649), (18509,-0.896426), (18510,-1.046404), (18511,-1.116483), (18512,-1.263204), (18513,-0.989561), (18514,-1.138143), (18515,-0.829197), (18516,-0.966169), (18517,-0.801680), (18518,-0.979059), (18519,-0.939521), (18520,-1.283654), (18521,-1.017907), (18522,-1.154410), (18523,-0.839427), (18524,-0.998228), (18525,-0.967976), (18526,-1.099376), (18527,-1.177814), (18528,-1.319896), (18529,-1.064368), (18530,-1.255216), (18531,-0.860341), (18532,-1.028427), (18533,-0.877876), (18534,-1.031567), (18535,-0.994816), (18536,-1.342199), (18537,-1.040686), (18538,-0.808846), (18539,-0.851523), (18540,-1.029835), (18541,-1.019095), (18542,-1.190438), (18543,-1.235432), (18544,-1.404452), (18545,-1.134529), (18546,-0.879464), (18547,-0.935141), (18548,-1.114849), (18549,-0.960579), (18550,-1.029268), (18551,-1.077049), (18552,-1.254898), (18553,-0.995187), (18554,-1.138196), (18555,-0.821817), (18556,-0.958789), (18557,-0.934573), (18558,-1.068296), (18559,-1.167172), (18560,-1.514562), (18561,-1.240913), (18562,-0.986318), (18563,-1.049897), (18564,-1.180827), (18565,-1.069293), (18566,-1.104532), (18567,-1.149996), (18568,-1.432352), (18569,-1.145703), (18570,-0.927332), (18571,-0.975120), (18572,-1.118128), (18573,-1.104138), (18574,-1.250860), (18575,-1.338127), (18576,-1.527122), (18577,-1.217249), (18578,-0.944996), (18579,-1.029940), (18580,-1.220794), (18581,-1.051658), (18582,-1.109665), (18583,-1.172311), (18584,-1.324149), (18585,-1.474584), (18586,-0.792185), (18587,-0.949595), (18588,-1.006669), (18589,-1.166866), (18590,-1.189569), (18591,-1.322822), (18592,-1.369213), (18593,-1.512222), (18594,-0.851651), (18595,-1.010915), (18596,-1.085177), (18597,-1.229582), (18598,-1.007961), (18599,-1.136568), (18600,-1.489524), (18601,-1.261867), (18602,-1.004949), (18603,-1.153061), (18604,-1.235218), (18605,-1.418640), (18606,-1.367023), (18607,-1.531860), (18608,-1.596836), (18609,-1.365459), (18610,-1.098785), (18611,-1.237611), (18612,-1.280289), (18613,-1.381489), (18614,-1.222115), (18615,-1.361868), (18616,-1.421734), (18617,-1.560096), (18618,-0.905562), (18619,-1.029066), (18620,-1.080566), (18621,-1.236117), (18622,-1.253711), (18623,-1.394860), (18624,-1.455653), (18625,-1.625599), (18626,-0.948310), (18627,-1.101068), (18628,-1.166507), (18629,-1.312302), (18630,-1.077212), (18631,-1.221147), (18632,-1.322347), (18633,-1.483471), (18634,-0.810364), (18635,-0.962196), (18636,-1.036457), (18637,-1.168320), (18638,-1.190560), (18639,-1.293619), (18640,-1.377167), (18641,-1.552229), (18642,-0.863325), (18643,-1.000760), (18644,-1.114965), (18645,-1.211525), (18646,-0.946241), (18647,-1.115261), (18648,-1.325620), (18649,-1.489067), (18650,-0.804345), (18651,-0.960359), (18652,-1.014183), (18653,-1.146973), (18654,-1.187328), (18655,-1.290850), (18656,-1.363722), (18657,-1.533668), (18658,-0.855452), (18659,-1.024002), (18660,-1.076899), (18661,-1.206902), (18662,-0.977385), (18663,-1.151978), (18664,-1.197906), (18665,-1.341841), (18666,-0.680344), (18667,-0.821493), (18668,-0.888792), (18669,-1.057342), (18670,-1.079118), (18671,-1.240242), (18672,-1.316827), (18673,-1.440787), (18674,-0.782546), (18675,-0.939024), (18676,-1.010036), (18677,-1.146538), (18678,-0.905876), (18679,-1.062816), (18680,-1.258774), (18681,-1.382741), (18682,-0.740285), (18683,-0.857283), (18684,-0.912497), (18685,-1.085236), (18686,-1.066136), (18687,-1.235149), (18688,-1.247640), (18689,-1.410617), (18690,-0.750053), (18691,-0.871227), (18692,-0.944092), (18693,-1.062017), (18694,-0.859907), (18695,-0.987124), (18696,-1.275979), (18697,-1.413415), (18698,-0.744485), (18699,-0.900036), (18700,-0.953860), (18701,-1.099192), (18702,-1.090305), (18703,-1.244929), (18704,-1.312685), (18705,-1.480778), (18706,-0.773294), (18707,-0.927449), (18708,-0.975700), (18709,-1.157262), (18710,-0.916129), (18711,-1.066107), (18712,-1.202146), (18713,-0.925717), (18714,-1.089627), (18715,-0.759316), (18716,-0.888850), (18717,-0.877646), (18718,-1.015545), (18719,-1.071228), (18720,-1.251857), (18721,-0.987506), (18722,-1.128655), (18723,-0.799734), (18724,-0.962248), (18725,-0.847927), (18726,-0.980253), (18727,-0.932820), (18728,-1.254192), (18729,-0.976830), (18730,-0.752422), (18731,-0.787204), (18732,-0.952041), (18733,-0.946410), (18734,-1.099174), (18735,-1.181795), (18736,-1.319695), (18737,-1.028863), (18738,-0.772872), (18739,-0.830878), (18740,-1.025909), (18741,-0.852127), (18742,-0.891092), (18743,-0.946775), (18744,-1.308091), (18745,-1.029338), (18746,-0.771951), (18747,-0.841573), (18748,-0.992941), (18749,-0.981730), (18750,-1.215784), (18751,-1.276577), (18752,-1.476717), (18753,-1.160338), (18754,-0.924779), (18755,-0.969316), (18756,-1.135549), (18757,-0.995681), (18758,-1.067619), (18759,-1.171605), (18760,-1.429347), (18761,-1.111578), (18762,-0.867659), (18763,-0.921946), (18764,-1.045913), (18765,-1.025417), (18766,-1.173535), (18767,-1.249656), (18768,-1.391732), (18769,-1.124589), (18770,-0.909473), (18771,-0.940073), (18772,-1.124884), (18773,-0.965504), (18774,-1.046272), (18775,-1.081054), (18776,-1.186436), (18777,-0.916970), (18778,-1.051156), (18779,-0.720844), (18780,-0.861993), (18781,-0.843820), (18782,-1.011444), (18783,-1.118686), (18784,-1.235220), (18785,-0.961107), (18786,-1.083215), (18787,-0.738502), (18788,-0.902412), (18789,-0.761616), (18790,-0.902765), (18791,-0.877160), (18792,-1.397334), (18793,-0.733050), (18794,-0.875132), (18795,-0.932206), (18796,-1.138388), (18797,-1.121142), (18798,-1.281802), (18799,-1.346772), (18800,-1.464696), (18801,-0.815741), (18802,-0.967109), (18803,-1.046480), (18804,-1.193209), (18805,-0.986916), (18806,-1.107627), (18807,-1.147049), (18808,-1.329537), (18809,-1.063327), (18810,-0.835206), (18811,-0.876951), (18812,-1.057586), (18813,-1.023152), (18814,-1.214006), (18815,-1.263647), (18816,-1.505126), (18817,-1.192930), (18818,-0.952267), (18819,-1.013060), (18820,-1.155136), (18821,-1.008298), (18822,-1.115540), (18823,-1.147536), (18824,-1.416423), (18825,-1.150676), (18826,-0.873777), (18827,-0.945252), (18828,-1.102662), (18829,-1.107714), (18830,-1.288343), (18831,-1.308259), (18832,-1.472633), (18833,-1.204099), (18834,-0.958791), (18835,-1.072069), (18836,-1.214614), (18837,-1.072886), (18838,-1.157367), (18839,-1.213513), (18840,-1.455926), (18841,-1.192032), (18842,-0.936968), (18843,-0.981042), (18844,-1.173286), (18845,-1.145358), (18846,-1.273038), (18847,-1.344513), (18848,-1.539544), (18849,-1.259858), (18850,-0.996434), (18851,-1.041899), (18852,-1.210918), (18853,-1.058044), (18854,-1.109545), (18855,-1.157332), (18856,-1.488924), (18857,-1.221317), (18858,-0.956960), (18859,-1.124589), (18860,-1.147293), (18861,-1.335817), (18862,-1.316254), (18863,-1.475518), (18864,-1.526092), (18865,-1.290076), (18866,-0.971373), (18867,-1.161295), (18868,-1.205363), (18869,-1.290776), (18870,-1.132323), (18871,-1.286478), (18872,-1.485228), (18873,-1.213908), (18874,-0.977885), (18875,-1.033568), (18876,-1.156602), (18877,-1.147721), (18878,-1.357148), (18879,-1.423050), (18880,-1.540975), (18881,-1.269191), (18882,-1.034565), (18883,-1.103254), (18884,-1.282956), (18885,-1.131935), (18886,-1.189941), (18887,-1.259557), (18888,-1.339861), (18889,-1.488443), (18890,-0.814404), (18891,-0.948583), (18892,-0.982438), (18893,-1.131483), (18894,-1.151400), (18895,-1.306018), (18896,-1.348232), (18897,-1.501460), (18898,-0.822311), (18899,-0.979252), (18900,-1.015424), (18901,-1.185377), (18902,-0.954927), (18903,-1.133702), (18904,-1.430460), (18905,-1.183291), (18906,-0.965383), (18907,-0.991343), (18908,-1.137601), (18909,-1.139866), (18910,-1.327928), (18911,-1.332052), (18912,-1.505718), (18913,-1.187016), (18914,-0.959822), (18915,-1.002964), (18916,-1.141789), (18917,-0.995878), (18918,-1.060854), (18919,-1.115141), (18920,-1.194512), (18921,-1.349136), (18922,-0.658835), (18923,-0.808813), (18924,-0.867747), (18925,-1.046985), (18926,-1.077121), (18927,-1.202478), (18928,-1.251192), (18929,-1.425785), (18930,-0.761038), (18931,-0.924021), (18932,-0.980631), (18933,-1.161723), (18934,-0.949858), (18935,-1.072892), (18936,-1.374759), (18937,-1.092287), (18938,-0.853948), (18939,-0.882687), (18940,-1.022909), (18941,-1.000090), (18942,-1.167256), (18943,-1.254524), (18944,-1.403569), (18945,-1.120170), (18946,-0.865105), (18947,-0.953769), (18948,-1.086552), (18949,-0.944360), (18950,-1.015836), (18951,-1.072916), (18952,-1.306499), (18953,-1.430460), (18954,-0.767109), (18955,-0.890607), (18956,-0.952326), (18957,-1.125529), (18958,-1.143122), (18959,-1.290308), (18960,-1.319517), (18961,-1.469025), (18962,-0.809851), (18963,-0.964932), (18964,-1.032231), (18965,-1.175239), (18966,-0.939680), (18967,-1.096621), (18968,-1.246135), (18969,-0.974815), (18970,-1.096453), (18971,-0.781934), (18972,-0.931442), (18973,-0.946249), (18974,-1.116202), (18975,-1.167702), (18976,-1.296309), (18977,-1.039855), (18978,-1.200045), (18979,-0.853942), (18980,-0.996018), (18981,-0.878447), (18982,-1.027029), (18983,-0.941968), (18984,-1.309790), (18985,-1.012459), (18986,-0.736493), (18987,-0.789384), (18988,-0.941221), (18989,-0.945809), (18990,-1.139444), (18991,-1.198840), (18992,-1.364147), (18993,-1.072852), (18994,-0.797349), (18995,-0.846063), (18996,-1.036918), (18997,-0.855703), (18998,-0.923002), (18999,-0.994014), (19000,-1.387383), (19001,-1.105838), (19002,-0.869821), (19003,-0.954302), (19004,-1.090805), (19005,-1.086107), (19006,-1.244438), (19007,-1.285262), (19008,-1.450563), (19009,-1.165304), (19010,-0.944616), (19011,-0.991470), (19012,-1.140515), (19013,-0.981142), (19014,-1.032179), (19015,-1.117586), (19016,-1.396693), (19017,-1.120263), (19018,-0.887490), (19019,-0.923199), (19020,-1.082463), (19021,-1.032242), (19022,-1.203585), (19023,-1.262518), (19024,-1.418996), (19025,-1.138847), (19026,-0.900044), (19027,-0.984525), (19028,-1.109418), (19029,-0.971403), (19030,-1.014081), (19031,-1.002877), (19032,-1.158892), (19033,-0.889425), (19034,-1.042653), (19035,-0.730457), (19036,-0.859990), (19037,-0.864115), (19038,-1.016416), (19039,-1.093928), (19040,-1.262947), (19041,-0.989768), (19042,-1.156001), (19043,-0.824757), (19044,-0.933395), (19045,-0.779588), (19046,-0.943498), (19047,-0.956915), (19048,-1.449219), (19049,-0.745455), (19050,-0.910755), (19051,-0.944141), (19052,-1.088546), (19053,-1.088951), (19054,-1.247752), (19055,-1.311795), (19056,-1.464559), (19057,-0.795166), (19058,-0.977654), (19059,-1.024509), (19060,-1.184242), (19061,-0.945896), (19062,-1.102844), (19063,-1.133443), (19064,-1.294566), (19065,-1.014417), (19066,-0.790010), (19067,-0.845224), (19068,-1.017030), (19069,-1.002576), (19070,-1.188321), (19071,-1.221706), (19072,-1.661061), (19073,-0.981449), (19074,-1.141640), (19075,-1.228444), (19076,-1.393280), (19077,-1.141009), (19078,-1.281694), (19079,-1.355486), (19080,-1.502678), (19081,-1.255046), (19082,-1.002768), (19083,-1.139270), (19084,-1.164297), (19085,-1.344462), (19086,-1.353233), (19087,-1.464658), (19088,-1.517548), (19089,-1.283855), (19090,-1.036223), (19091,-1.198273), (19092,-1.241878), (19093,-1.305921), (19094,-1.140041), (19095,-1.305811), (19096,-1.321545), (19097,-1.503107), (19098,-0.829067), (19099,-0.999014), (19100,-1.051447), (19101,-1.206992), (19102,-1.184642), (19103,-1.353199), (19104,-1.387511), (19105,-1.540275), (19106,-0.839761), (19107,-0.994379), (19108,-1.072360), (19109,-1.210260), (19110,-0.984456), (19111,-1.121892), (19112,-1.348969), (19113,-1.083222), (19114,-0.813756), (19115,-0.978599), (19116,-1.046355), (19117,-1.187974), (19118,-1.197671), (19119,-1.375977), (19120,-1.435373), (19121,-1.197961), (19122,-0.937323), (19123,-1.087301), (19124,-1.123473), (19125,-1.202381), (19126,-1.031392), (19127,-1.177650), (19128,-1.508315), (19129,-1.261610), (19130,-0.983784), (19131,-1.153267), (19132,-1.220566), (19133,-1.443461), (19134,-1.432257), (19135,-1.545072), (19136,-1.616547), (19137,-1.362416), (19138,-1.068798), (19139,-1.229922), (19140,-1.323225), (19141,-1.382158), (19142,-1.215352), (19143,-1.351855), (19144,-1.442372), (19145,-1.204959), (19146,-0.941071), (19147,-1.071538), (19148,-1.144403), (19149,-1.333861), (19150,-1.317085), (19151,-1.484708), (19152,-1.542251), (19153,-1.311807), (19154,-1.060919), (19155,-1.200215), (19156,-1.214089), (19157,-1.271169), (19158,-1.142446), (19159,-1.286844), (19160,-1.343924), (19161,-1.525016), (19162,-0.832399), (19163,-0.974481), (19164,-1.033414), (19165,-1.165734), (19166,-1.187510), (19167,-1.346774), (19168,-1.404781), (19169,-1.555685), (19170,-0.881646), (19171,-1.026978), (19172,-1.104489), (19173,-1.246571), (19174,-1.010548), (19175,-1.145661), (19176,-1.212490), (19177,-1.355036), (19178,-0.683319), (19179,-0.829578), (19180,-0.901053), (19181,-1.035696), (19182,-1.032388), (19183,-1.197231), (19184,-1.261737), (19185,-1.415892), (19186,-0.747889), (19187,-0.914592), (19188,-0.985134), (19189,-1.128143), (19190,-0.856823), (19191,-1.010044), (19192,-1.117756), (19193,-1.290489), (19194,-0.619236), (19195,-0.769677), (19196,-0.817464), (19197,-0.999026), (19198,-1.015223), (19199,-1.209327), (19200,-1.213916), (19201,-1.365284), (19202,-0.711682), (19203,-0.859800), (19204,-0.936385), (19205,-1.084967), (19206,-0.847554), (19207,-0.959899), (19208,-1.191629), (19209,-1.378301), (19210,-0.701475), (19211,-0.851910), (19212,-0.892728), (19213,-1.014835), (19214,-1.048691), (19215,-1.185193), (19216,-1.222762), (19217,-1.362514), (19218,-0.712632), (19219,-0.873287), (19220,-0.941512), (19221,-1.096130), (19222,-0.879155), (19223,-1.028670), (19224,-1.404387), (19225,-1.120988), (19226,-0.880789), (19227,-0.943905), (19228,-1.054397), (19229,-1.034827), (19230,-1.217322), (19231,-1.272999), (19232,-1.432733), (19233,-1.184168), (19234,-0.899842), (19235,-0.952739), (19236,-1.123149), (19237,-0.963306), (19238,-1.022709), (19239,-1.087678), (19240,-1.300360), (19241,-0.996524), (19242,-0.746105), (19243,-0.813867), (19244,-1.000996), (19245,-0.960994), (19246,-1.189469), (19247,-1.251658), (19248,-1.391411), (19249,-1.095006), (19250,-0.831582), (19251,-0.877973), (19252,-1.091582), (19253,-0.984694), (19254,-1.061279), (19255,-1.114176), (19256,-1.361692), (19257,-1.029991), (19258,-0.779103), (19259,-0.846401), (19260,-1.033536), (19261,-0.993529), (19262,-1.186236), (19263,-1.247029), (19264,-1.432774), (19265,-1.133113), (19266,-0.878049), (19267,-0.943488), (19268,-1.097642), (19269,-0.908075), (19270,-0.959112), (19271,-1.018509), (19272,-1.295292), (19273,-0.990991), (19274,-0.739640), (19275,-0.795323), (19276,-1.010329), (19277,-0.984260), (19278,-1.148170), (19279,-1.213609), (19280,-1.383092), (19281,-1.125241), (19282,-0.870176), (19283,-0.899379), (19284,-1.059576), (19285,-0.907629), (19286,-0.985140), (19287,-1.058012), (19288,-1.400749), (19289,-1.104345), (19290,-0.869255), (19291,-0.944913), (19292,-1.093495), (19293,-1.052097), (19294,-1.203465), (19295,-1.248930), (19296,-1.421662), (19297,-1.126655), (19298,-0.880413), (19299,-0.929127), (19300,-1.092574), (19301,-0.954101), (19302,-1.048331), (19303,-1.097515), (19304,-1.390090), (19305,-0.693753), (19306,-0.800532), (19307,-0.841350), (19308,-0.968567), (19309,-1.017281), (19310,-1.192337), (19311,-1.219223), (19312,-1.385919), (19313,-0.691442), (19314,-0.859998), (19315,-0.918005), (19316,-1.068439), (19317,-0.869116), (19318,-1.023734), (19319,-1.058053), (19320,-1.480683), (19321,-0.804326), (19322,-0.960804), (19323,-1.022060), (19324,-1.174355), (19325,-1.195668), (19326,-1.369797), (19327,-1.446382), (19328,-1.486737), (19329,-1.631136), (19330,-0.952913), (19331,-1.109861), (19332,-1.181336), (19333,-1.327131), (19334,-1.085999), (19335,-1.214142), (19336,-1.378052), (19337,-1.509915), (19338,-0.854454), (19339,-0.974238), (19340,-1.048500), (19341,-1.209624), (19342,-1.252765), (19343,-1.385548), (19344,-1.449597), (19345,-1.603752), (19346,-0.934822), (19347,-1.078757), (19348,-1.142337), (19349,-1.297888), (19350,-1.071620), (19351,-1.235067), (19352,-1.471437), (19353,-1.494140), (19354,-1.245575), (19355,-0.939885), (19356,-1.093576), (19357,-1.142754), (19358,-1.341967), (19359,-1.328440), (19360,-1.466803), (19361,-1.498329), (19362,-1.314334), (19363,-1.073202), (19364,-1.224570), (19365,-1.265394), (19366,-1.314572), (19367,-1.146369), (19368,-1.356728), (19369,-1.421698), (19370,-1.194040), (19371,-0.903209), (19372,-1.043895), (19373,-1.084713), (19374,-1.305291), (19375,-1.289905), (19376,-1.455211), (19377,-1.494633), (19378,-1.237245), (19379,-0.948274), (19380,-1.121013), (19381,-1.163221), (19382,-1.203576), (19383,-1.060921), (19384,-1.400408), (19385,-1.459805), (19386,-1.215892), (19387,-0.951535), (19388,-1.121018), (19389,-1.150691), (19390,-1.301595), (19391,-1.277386), (19392,-1.466380), (19393,-1.490010), (19394,-1.274895), (19395,-1.017044), (19396,-1.190704), (19397,-1.263575), (19398,-1.331331), (19399,-1.150123), (19400,-1.346550), (19401,-1.414769), (19402,-1.175966), (19403,-0.896281), (19404,-1.043009), (19405,-1.065242), (19406,-1.227299), (19407,-1.220272), (19408,-1.385109), (19409,-1.425000), (19410,-1.208952), (19411,-0.932986), (19412,-1.087610), (19413,-1.185560), (19414,-1.243566), (19415,-1.084186), (19416,-1.503103), (19417,-1.576438), (19418,-1.332056), (19419,-1.045870), (19420,-1.201421), (19421,-1.238983), (19422,-1.437270), (19423,-1.420487), (19424,-1.551423), (19425,-1.602924), (19426,-1.353895), (19427,-1.089075), (19428,-1.238126), (19429,-1.323534), (19430,-1.357853), (19431,-1.241202), (19432,-1.342871), (19433,-1.411097), (19434,-1.186689), (19435,-0.895395), (19436,-1.024934), (19437,-1.065283), (19438,-1.246845), (19439,-1.242610), (19440,-1.406057), (19441,-1.428760), (19442,-1.223394), (19443,-0.912588), (19444,-1.070462), (19445,-1.114994), (19446,-1.174860), (19447,-1.068898), (19448,-1.111113), (19449,-1.169113), (19450,-1.332560), (19451,-0.707292), (19452,-0.836369), (19453,-0.886473), (19454,-1.040634), (19455,-1.068447), (19456,-1.183115), (19457,-1.218824), (19458,-1.364155), (19459,-0.687329), (19460,-0.821515), (19461,-0.872089), (19462,-1.014628), (19463,-0.795794), (19464,-1.142714), (19465,-1.212336), (19466,-1.326077), (19467,-0.684091), (19468,-0.855898), (19469,-0.938982), (19470,-1.053193), (19471,-1.090762), (19472,-1.256062), (19473,-1.297813), (19474,-1.413414), (19475,-0.750057), (19476,-0.917217), (19477,-0.971041), (19478,-1.114050), (19479,-0.886856), (19480,-1.152023), (19481,-1.327086), (19482,-1.032535), (19483,-0.774684), (19484,-0.802496), (19485,-0.955261), (19486,-0.959849), (19487,-1.134905), (19488,-1.193838), (19489,-1.370754), (19490,-1.085502), (19491,-0.814182), (19492,-0.937216), (19493,-1.064889), (19494,-0.886931), (19495,-0.947261), (19496,-1.260274), (19497,-1.424184), (19498,-0.768259), (19499,-0.912664), (19500,-0.968342), (19501,-1.126215), (19502,-1.140559), (19503,-1.336053), (19504,-1.400096), (19505,-1.536135), (19506,-0.865352), (19507,-1.020897), (19508,-1.097482), (19509,-1.186609), (19510,-0.965921), (19511,-1.141440), (19512,-1.151137), (19513,-1.338735), (19514,-1.019107), (19515,-0.778907), (19516,-0.850383), (19517,-1.012433), (19518,-0.985901), (19519,-1.154920), (19520,-1.208744), (19521,-1.339211), (19522,-1.084146), (19523,-0.843020), (19524,-0.893124), (19525,-1.036133), (19526,-0.879545), (19527,-0.956130), (19528,-1.106102), (19529,-1.283944), (19530,-1.014947), (19531,-0.764066), (19532,-0.799774), (19533,-0.960898), (19534,-0.958054), (19535,-1.132646), (19536,-1.173464), (19537,-1.324369), (19538,-1.058622), (19539,-0.826782), (19540,-0.872246), (19541,-1.019895), (19542,-0.874917), (19543,-0.942679), (19544,-1.084291), (19545,-1.234732), (19546,-0.959230), (19547,-0.726926), (19548,-0.783536), (19549,-0.920972), (19550,-0.912555), (19551,-1.107585), (19552,-1.140971), (19553,-1.285370), (19554,-1.029842), (19555,-0.804508), (19556,-0.845789), (19557,-0.981828), (19558,-0.827095), (19559,-0.921331), (19560,-1.204614), (19561,-1.329971), (19562,-0.654541), (19563,-0.781288), (19564,-0.875525), (19565,-1.020393), (19566,-1.031018), (19567,-1.191678), (19568,-1.226923), (19569,-1.366213), (19570,-0.686600), (19571,-0.826823), (19572,-0.890402), (19573,-1.063135), (19574,-0.853129), (19575,-1.004961), (19576,-1.277561), (19577,-1.420106), (19578,-0.723769), (19579,-0.887216), (19580,-0.957295), (19581,-1.115168), (19582,-1.142981), (19583,-1.287850), (19584,-1.628264), (19585,-1.782888), (19586,-1.095373), (19587,-1.238382), (19588,-1.341911), (19589,-1.504888), (19590,-1.270261), (19591,-1.420703), (19592,-1.498684), (19593,-1.639363), (19594,-0.947678), (19595,-1.091614), (19596,-1.148687), (19597,-1.300055), (19598,-1.309290), (19599,-1.484352), (19600,-1.546535), (19601,-1.693257), (19602,-1.003425), (19603,-1.159903), (19604,-1.216983), (19605,-1.349303), (19606,-1.095634), (19607,-1.267904), (19608,-1.482446), (19609,-1.526514), (19610,-1.291887), (19611,-1.009415), (19612,-1.180295), (19613,-1.227155), (19614,-1.413357), (19615,-1.385435), (19616,-1.546552), (19617,-1.623607), (19618,-1.396876), (19619,-1.086070), (19620,-1.208641), (19621,-1.292658), (19622,-1.394791), (19623,-1.240057), (19624,-1.460635), (19625,-1.478692), (19626,-1.267290), (19627,-0.969489), (19628,-1.152448), (19629,-1.177937), (19630,-1.371108), (19631,-1.360368), (19632,-1.489908), (19633,-1.548377), (19634,-1.299349), (19635,-1.019670), (19636,-1.217023), (19637,-1.276420), (19638,-1.284721), (19639,-1.096544), (19640,-1.544264), (19641,-1.611557), (19642,-1.353706), (19643,-1.083313), (19644,-1.228644), (19645,-1.288041), (19646,-1.486791), (19647,-1.423559), (19648,-1.610230), (19649,-1.645939), (19650,-1.403880), (19651,-1.111658), (19652,-1.281605), (19653,-1.378628), (19654,-1.452426), (19655,-1.267035), (19656,-1.394715), (19657,-1.467587), (19658,-1.221808), (19659,-0.936087), (19660,-1.101393), (19661,-1.131529), (19662,-1.312158), (19663,-1.285625), (19664,-1.428171), (19665,-1.487567), (19666,-1.234826), (19667,-0.946317), (19668,-1.120447), (19669,-1.204927), (19670,-1.245282), (19671,-1.087762), (19672,-1.456980), (19673,-1.542387), (19674,-1.304511), (19675,-1.016003), (19676,-1.150652), (19677,-1.228627), (19678,-1.399970), (19679,-1.390156), (19680,-1.570328), (19681,-1.623688), (19682,-1.360258), (19683,-1.073146), (19684,-1.215691), (19685,-1.309922), (19686,-1.368861), (19687,-1.217840), (19688,-1.358063), (19689,-1.421179), (19690,-1.171224), (19691,-0.868313), (19692,-1.035010), (19693,-1.086511), (19694,-1.254140), (19695,-1.252222), (19696,-1.402200), (19697,-1.517338), (19698,-1.261341), (19699,-0.978875), (19700,-1.145108), (19701,-1.212864), (19702,-1.265298), (19703,-1.124959), (19704,-1.152772), (19705,-1.200560), (19706,-1.337069), (19707,-0.681608), (19708,-0.859450), (19709,-0.924889), (19710,-1.067434), (19711,-1.059944), (19712,-1.223854), (19713,-1.277678), (19714,-1.422076), (19715,-0.730855), (19716,-0.904521), (19717,-0.998751), (19718,-1.147333), (19719,-0.893201), (19720,-1.248480), (19721,-1.280476), (19722,-1.431844), (19723,-0.761987), (19724,-0.924964), (19725,-0.974148), (19726,-1.138522), (19727,-1.157042), (19728,-1.284722), (19729,-1.310675), (19730,-1.453684), (19731,-0.786150), (19732,-0.955170), (19733,-1.031755), (19734,-1.227712), (19735,-0.962892), (19736,-1.230852), (19737,-1.414267), (19738,-1.122046), (19739,-0.921326), (19740,-0.949139), (19741,-1.094471), (19742,-1.087444), (19743,-1.235562), (19744,-1.289385), (19745,-1.467698), (19746,-1.201481), (19747,-0.997981), (19748,-1.050872), (19749,-1.166010), (19750,-1.005703), (19751,-1.106445), (19752,-1.392051), (19753,-1.568967), (19754,-0.874953), (19755,-1.028644), (19756,-1.088510), (19757,-1.223616), (19758,-1.226814), (19759,-1.376786), (19760,-1.438512), (19761,-1.560150), (19762,-0.866142), (19763,-1.004504), (19764,-1.074583), (19765,-1.221305), (19766,-0.998294), (19767,-1.171960), (19768,-1.218814), (19769,-1.335349), (19770,-1.074241), (19771,-0.838225), (19772,-0.856282), (19773,-1.014156), (19774,-0.980654), (19775,-1.194263), (19776,-1.234155), (19777,-1.405028), (19778,-1.111410), (19779,-0.901404), (19780,-0.978452), (19781,-1.115425), (19782,-0.963014), (19783,-1.052604), (19784,-1.175638), (19785,-1.334439), (19786,-1.058473), (19787,-0.831273), (19788,-0.900895), (19789,-1.081060), (19790,-1.048491), (19791,-1.206822), (19792,-1.273658), (19793,-1.425026), (19794,-1.132335), (19795,-0.890739), (19796,-0.947819), (19797,-1.099650), (19798,-0.948166), (19799,-1.012679), (19800,-1.210496), (19801,-1.408776), (19802,-1.112372), (19803,-0.854521), (19804,-0.895339), (19805,-1.072718), (19806,-1.061051), (19807,-1.198487), (19808,-1.283894), (19809,-1.443621), (19810,-1.169978), (19811,-0.941388), (19812,-0.991035), (19813,-1.120105), (19814,-0.972341), (19815,-1.047999), (19816,-1.329422), (19817,-1.535605), (19818,-0.835091), (19819,-0.982739), (19820,-1.017985), (19821,-1.159603), (19822,-1.166508), (19823,-1.313700), (19824,-1.414436), (19825,-1.570450), (19826,-0.883869), (19827,-0.975782), (19828,-1.046331), (19829,-1.205131), (19830,-1.006735), (19831,-1.124196), (19832,-1.437672), (19833,-1.592760), (19834,-0.927543), (19835,-1.068229), (19836,-1.140167), (19837,-1.316620), (19838,-1.338859), (19839,-1.467003), (19840,-1.512004), (19841,-1.676377), (19842,-1.405051), (19843,-1.143024), (19844,-1.194524), (19845,-1.344502), (19846,-1.196268), (19847,-1.244055), (19848,-1.435836), (19849,-1.603459), (19850,-1.311238), (19851,-1.082648), (19852,-1.138794), (19853,-1.289236), (19854,-1.297074), (19855,-1.460984), (19856,-1.559403), (19857,-1.710771), (19858,-1.419940), (19859,-1.185313), (19860,-1.237277), (19861,-1.383072), (19862,-1.239484), (19863,-1.287272), (19864,-1.434000), (19865,-1.484567), (19866,-1.646154), (19867,-0.950287), (19868,-1.101192), (19869,-1.155479), (19870,-1.292451), (19871,-1.303539), (19872,-1.464199), (19873,-1.529638), (19874,-1.688439), (19875,-1.021832), (19876,-1.165304), (19877,-1.201013), (19878,-1.362136), (19879,-1.125650), (19880,-1.566395), (19881,-1.641590), (19882,-1.371197), (19883,-1.110096), (19884,-1.258677), (19885,-1.319934), (19886,-1.468515), (19887,-1.444306), (19888,-1.623538), (19889,-1.674576), (19890,-1.433449), (19891,-1.199286), (19892,-1.372025), (19893,-1.428172), (19894,-1.516830), (19895,-1.363492), (19896,-1.526939), (19897,-1.605377), (19898,-1.763251), (19899,-1.071097), (19900,-1.198313), (19901,-1.250277), (19902,-1.427656), (19903,-1.392301), (19904,-1.510689), (19905,-1.597956), (19906,-1.755830), (19907,-1.087364), (19908,-1.252670), (19909,-1.300921), (19910,-1.471331), (19911,-1.243673), (19912,-1.407584), (19913,-1.462797), (19914,-1.598837), (19915,-0.921547), (19916,-1.043191), (19917,-1.114667), (19918,-1.270218), (19919,-1.278982), (19920,-1.415955), (19921,-1.470705), (19922,-1.657376), (19923,-0.989373), (19924,-1.133778), (19925,-1.176919), (19926,-1.338507), (19927,-1.077406), (19928,-1.406674), (19929,-1.464211), (19930,-1.617902), (19931,-0.949905), (19932,-1.099413), (19933,-1.129086), (19934,-1.279990), (19935,-1.285042), (19936,-1.472640), (19937,-1.522287), (19938,-1.677368), (19939,-0.988933), (19940,-1.122650), (19941,-1.218276), (19942,-1.384973), (19943,-1.128982), (19944,-1.278959), (19945,-1.364830), (19946,-1.487401), (19947,-0.787351), (19948,-0.936395), (19949,-0.983256), (19950,-1.148093), (19951,-1.164760), (19952,-1.329597), (19953,-1.373665), (19954,-1.562659), (19955,-0.882584), (19956,-1.026519), (19957,-1.065014), (19958,-1.209419), (19959,-0.989188), (19960,-1.280836), (19961,-1.326764), (19962,-1.469309), (19963,-0.835213), (19964,-0.995410), (19965,-1.013004), (19966,-1.176914), (19967,-1.202867), (19968,-1.305463), (19969,-1.361610), (19970,-1.521807), (19971,-0.845907), (19972,-0.990306), (19973,-1.046459), (19974,-1.188072), (19975,-0.959945), (19976,-1.291536), (19977,-1.350939), (19978,-1.516702), (19979,-0.812012), (19980,-0.956411), (19981,-1.047861), (19982,-1.189473), (19983,-1.235864), (19984,-1.394665), (19985,-1.457318), (19986,-1.609149), (19987,-0.948115), (19988,-1.108775), (19989,-1.151917), (19990,-1.289353), (19991,-1.063549), (19992,-1.340795), (19993,-1.529790), (19994,-1.216197), (19995,-0.969492), (19996,-1.005670), (19997,-1.168184), (19998,-1.180668), (19999,-1.342255), (20000,-1.367281), (20001,-1.532588), (20002,-1.242220), (20003,-1.005734), (20004,-1.043765), (20005,-1.216504), (20006,-1.031113), (20007,-1.119771), (20008,-1.214940), (20009,-1.361662), (20010,-1.103811), (20011,-0.871508), (20012,-0.929514), (20013,-1.090168), (20014,-1.085470), (20015,-1.229406), (20016,-1.291589), (20017,-1.456425), (20018,-1.195325), (20019,-0.935150), (20020,-0.996870), (20021,-1.170536), (20022,-1.024168), (20023,-1.111898), (20024,-1.325044), (20025,-1.468979), (20026,-1.207878), (20027,-0.976502), (20028,-1.037758), (20029,-1.170084), (20030,-1.178386), (20031,-1.335326), (20032,-1.370572), (20033,-1.528446), (20034,-1.261772), (20035,-1.015530), (20036,-1.071213), (20037,-1.184955), (20038,-1.085963), (20039,-1.111452), (20040,-1.289301), (20041,-1.463893), (20042,-1.202323), (20043,-0.940759), (20044,-0.982040), (20045,-1.139914), (20046,-1.114772), (20047,-1.292151), (20048,-1.311141), (20049,-1.499666), (20050,-1.206517), (20051,-0.952843), (20052,-1.043366), (20053,-1.239324), (20054,-1.041390), (20055,-1.116585), (20056,-1.259124), (20057,-1.431394), (20058,-1.129880), (20059,-0.914765), (20060,-0.946297), (20061,-1.093019), (20062,-1.081815), (20063,-1.249902), (20064,-1.318591), (20065,-1.475531), (20066,-1.216290), (20067,-0.968658), (20068,-1.045243), (20069,-1.191965), (20070,-1.050237), (20071,-1.098487), (20072,-1.364588), (20073,-1.503877), (20074,-0.826588), (20075,-0.990498), (20076,-1.025280), (20077,-1.173392), (20078,-1.215143), (20079,-1.388339), (20080,-1.458425), (20081,-1.564270), (20082,-0.912065), (20083,-1.082475), (20084,-1.160920), (20085,-1.304855), (20086,-1.042364), (20087,-1.198372), (20088,-1.286572), (20089,-1.435617), (20090,-1.148505), (20091,-0.928274), (20092,-0.995573), (20093,-1.190604), (20094,-1.119013), (20095,-1.312183), (20096,-1.615441), (20097,-1.670661), (20098,-1.427212), (20099,-1.119655), (20100,-1.282176), (20101,-1.346218), (20102,-1.432559), (20103,-1.283861), (20104,-1.448698), (20105,-1.498809), (20106,-1.258146), (20107,-0.991929), (20108,-1.114500), (20109,-1.185048), (20110,-1.373110), (20111,-1.339614), (20112,-1.490513), (20113,-1.568031), (20114,-1.334794), (20115,-1.037000), (20116,-1.166997), (20117,-1.259380), (20118,-1.313204), (20119,-1.180761), (20120,-1.524431), (20121,-1.596370), (20122,-1.342702), (20123,-1.065339), (20124,-1.218567), (20125,-1.265428), (20126,-1.459525), (20127,-1.410232), (20128,-1.555100), (20129,-1.660946), (20130,-1.430966), (20131,-1.163359), (20132,-1.281753), (20133,-1.301200), (20134,-1.367566), (20135,-1.223984), (20136,-1.335866), (20137,-1.489094), (20138,-1.111407), (20139,-1.263701), (20140,-1.002601), (20141,-1.154432), (20142,-1.233803), (20143,-1.390744), (20144,-1.385583), (20145,-1.519299), (20146,-1.164367), (20147,-1.310626), (20148,-1.028623), (20149,-1.181381), (20150,-1.161818), (20151,-1.335484), (20152,-1.451549), (20153,-1.595484), (20154,-1.248448), (20155,-1.406322), (20156,-1.132216), (20157,-1.266395), (20158,-1.360169), (20159,-1.512927), (20160,-1.497077), (20161,-1.653554), (20162,-1.317670), (20163,-1.512237), (20164,-1.231625), (20165,-1.374634), (20166,-1.359247), (20167,-1.509689), (20168,-1.285744), (20169,-1.445472), (20170,-1.130026), (20171,-1.253060), (20172,-1.017037), (20173,-1.153546), (20174,-1.232917), (20175,-1.358274), (20176,-1.347997), (20177,-1.486360), (20178,-1.131428), (20179,-1.306484), (20180,-0.993361), (20181,-1.147979), (20182,-1.108904), (20183,-1.286283), (20184,-1.373087), (20185,-1.562081), (20186,-1.215978), (20187,-1.352481), (20188,-1.085338), (20189,-1.257144), (20190,-1.328619), (20191,-1.489279), (20192,-1.453924), (20193,-1.603433), (20194,-1.252683), (20195,-1.414271), (20196,-1.133195), (20197,-1.276667), (20198,-1.261280), (20199,-1.404289), (20200,-1.292285), (20201,-1.466884), (20202,-1.118451), (20203,-1.262856), (20204,-0.998499), (20205,-1.158696), (20206,-1.227849), (20207,-1.397332), (20208,-1.382408), (20209,-1.522167), (20210,-1.197429), (20211,-1.335328), (20212,-1.043100), (20213,-1.207474), (20214,-1.176295), (20215,-1.325810), (20216,-1.073995), (20217,-1.245801), (20218,-1.292656), (20219,-1.026909), (20220,-0.755125), (20221,-0.890701), (20222,-0.937092), (20223,-1.119581), (20224,-1.097231), (20225,-1.248136), (20226,-1.297777), (20227,-1.050608), (20228,-0.750028), (20229,-0.926010), (20230,-0.974724), (20231,-1.033194), (20232,-1.048934), (20233,-1.241642), (20234,-1.284320), (20235,-1.072918), (20236,-0.793696), (20237,-0.915803), (20238,-0.956621), (20239,-1.140506), (20240,-1.116297), (20241,-1.291353), (20242,-1.336354), (20243,-1.081752), (20244,-0.793244), (20245,-0.969696), (20246,-1.022593), (20247,-1.127043), (20248,-1.169720), (20249,-1.226331), (20250,-1.379095), (20251,-0.732463), (20252,-0.895910), (20253,-0.945551), (20254,-1.097852), (20255,-1.082928), (20256,-1.225937), (20257,-1.302985), (20258,-1.460859), (20259,-0.783564), (20260,-0.917750), (20261,-0.995261), (20262,-1.155922), (20263,-0.911076), (20264,-1.352291), (20265,-1.426552), (20266,-1.212364), (20267,-0.915496), (20268,-1.044103), (20269,-1.108146), (20270,-1.282275), (20271,-1.277108), (20272,-1.419183), (20273,-1.514353), (20274,-1.253246), (20275,-0.996791), (20276,-1.149086), (20277,-1.158783), (20278,-1.243734), (20279,-1.094109), (20280,-1.198559), (20281,-1.287686), (20282,-1.400501), (20283,-0.744582), (20284,-0.873189), (20285,-0.930726), (20286,-1.061656), (20287,-1.066714), (20288,-1.224118), (20289,-1.298843), (20290,-1.433029), (20291,-0.797080), (20292,-0.948448), (20293,-1.006917), (20294,-1.129951), (20295,-0.897178), (20296,-1.166065), (20297,-1.221285), (20298,-1.381476), (20299,-0.700937), (20300,-0.854628), (20301,-0.915884), (20302,-1.073758), (20303,-1.078347), (20304,-1.231105), (20305,-1.292824), (20306,-1.422364), (20307,-0.759477), (20308,-0.908985), (20309,-0.970705), (20310,-1.123006), (20311,-0.883733), (20312,-1.108024), (20313,-1.186469), (20314,-1.341550), (20315,-0.651255), (20316,-0.814702), (20317,-0.888501), (20318,-1.000852), (20319,-0.991971), (20320,-1.171204), (20321,-1.241752), (20322,-1.407986), (20323,-0.733946), (20324,-0.922941), (20325,-0.987447), (20326,-1.127206), (20327,-0.879574), (20328,-1.274796), (20329,-1.363460), (20330,-1.098640), (20331,-0.824070), (20332,-0.971255), (20333,-1.042267), (20334,-1.219646), (20335,-1.170352), (20336,-1.342628), (20337,-1.384836), (20338,-1.105157), (20339,-0.853806), (20340,-0.992632), (20341,-1.047388), (20342,-1.112827), (20343,-0.985495), (20344,-1.387229), (20345,-1.433620), (20346,-1.185055), (20347,-0.895620), (20348,-1.050238), (20349,-1.115214), (20350,-1.331146), (20351,-1.326912), (20352,-1.302233), (20353,-0.937088), (20354,-1.116320), (20355,-0.858939), (20356,-0.958748), (20357,-0.926637), (20358,-1.105875), (20359,-0.939996), (20360,-1.165220), (20361,-0.835372), (20362,-0.976985), (20363,-0.743285), (20364,-0.870965), (20365,-0.973097), (20366,-1.114246), (20367,-1.100720), (20368,-1.254411), (20369,-0.922240), (20370,-1.057816), (20371,-0.810184), (20372,-0.942973), (20373,-0.926660), (20374,-1.077101), (20375,-0.971140), (20376,-0.999416), (20377,-1.151711), (20378,-0.799102), (20379,-0.887302), (20380,-0.611799), (20381,-0.775709), (20382,-0.846258), (20383,-1.000876), (20384,-0.976666), (20385,-1.152649), (20386,-0.804686), (20387,-0.930507), (20388,-0.704709), (20389,-0.844462), (20390,-0.818862), (20391,-0.949792), (20392,-0.962276), (20393,-0.734149), (20394,-0.774504), (20395,-0.948633), (20396,-0.654552), (20397,-0.850510), (20398,-0.895511), (20399,-1.032013), (20400,-1.023133), (20401,-0.787116), (20402,-0.842330), (20403,-0.999277), (20404,-0.693581), (20405,-0.789677), (20406,-0.870901), (20407,-0.994405), (20408,-1.093745), (20409,-0.846582), (20410,-0.901333), (20411,-1.055024), (20412,-0.794386), (20413,-0.952724), (20414,-1.010724), (20415,-1.182067), (20416,-1.186655), (20417,-0.902329), (20418,-0.951043), (20419,-1.132605), (20420,-0.889619), (20421,-0.935084), (20422,-0.983335), (20423,-1.163963), (20424,-1.090982), (20425,-0.859605), (20426,-0.921794), (20427,-1.052255), (20428,-0.764216), (20429,-0.934163), (20430,-1.002388), (20431,-1.119379), (20432,-1.126291), (20433,-0.867513), (20434,-0.910654), (20435,-1.063882), (20436,-0.796738), (20437,-0.871464), (20438,-0.924824), (20439,-1.079911), (20440,-0.947939), (20441,-1.126244), (20442,-0.798720), (20443,-0.940802), (20444,-0.644861), (20445,-0.802728), (20446,-0.889532), (20447,-1.011176), (20448,-1.028770), (20449,-1.180138), (20450,-0.846107), (20451,-1.027669), (20452,-0.756813), (20453,-0.887279), (20454,-0.867716), (20455,-1.026047), (20456,-0.941456), (20457,-1.063094), (20458,-0.742075), (20459,-0.866962), (20460,-0.589606), (20461,-0.760479), (20462,-0.866795), (20463,-1.015840), (20464,-0.987448), (20465,-1.164363), (20466,-0.818723), (20467,-0.947800), (20468,-0.691339), (20469,-0.844567), (20470,-0.795273), (20471,-0.951287), (20472,-0.821168), (20473,-0.983688), (20474,-0.643158), (20475,-0.760613), (20476,-0.509268), (20477,-0.638338), (20478,-0.725142), (20479,-0.883016), (20480,-0.849051), (20481,-1.025040), (20482,-0.678003), (20483,-0.842840), (20484,-0.549686), (20485,-0.737754), (20486,-0.707038), (20487,-0.851907), (20488,-0.884829), (20489,-1.011113), (20490,-0.665936), (20491,-0.797793), (20492,-0.540412), (20493,-0.711748), (20494,-0.760469), (20495,-0.922982), (20496,-0.944289), (20497,-1.118888), (20498,-0.746768), (20499,-0.913001), (20500,-0.635638), (20501,-0.779110), (20502,-0.768370), (20503,-0.857497), (20504,-0.943374), (20505,-0.986515), (20506,-0.775577), (20507,-0.492641), (20508,-0.641223), (20509,-0.731277), (20510,-0.870572), (20511,-0.843576), (20512,-1.007950), (20513,-1.069670), (20514,-0.819715), (20515,-0.505659), (20516,-0.681648), (20517,-0.714570), (20518,-0.802300), (20519,-0.665218), (20520,-0.955933), (20521,-1.020440), (20522,-0.791856), (20523,-0.538181), (20524,-0.682123), (20525,-0.747092), (20526,-0.900320), (20527,-0.867745), (20528,-1.023759), (20529,-1.083162), (20530,-0.823915), (20531,-0.551198), (20532,-0.696993), (20533,-0.754073), (20534,-0.840407), (20535,-0.704258), (20536,-0.950384), (20537,-1.005135), (20538,-0.763075), (20539,-0.499651), (20540,-0.633368), (20541,-0.704843), (20542,-0.891514), (20543,-0.878914), (20544,-1.045147), (20545,-1.071570), (20546,-0.856912), (20547,-0.563294), (20548,-0.719308), (20549,-0.754554), (20550,-0.835321), (20551,-0.675015), (20552,-0.904879), (20553,-0.963349), (20554,-0.727332), (20555,-0.443934), (20556,-0.582759), (20557,-0.612432), (20558,-0.806999), (20559,-0.794399), (20560,-0.973638), (20561,-1.035357), (20562,-0.786799), (20563,-0.489461), (20564,-0.636183), (20565,-0.669575), (20566,-0.763805), (20567,-0.589103), (20568,-0.855197), (20569,-0.908094), (20570,-0.702735), (20571,-0.434665), (20572,-0.554443), (20573,-0.605949), (20574,-0.797261), (20575,-0.781411), (20576,-0.926279), (20577,-0.970347), (20578,-0.719002), (20579,-0.425847), (20580,-0.607873), (20581,-0.631039), (20582,-0.714130), (20583,-0.611881), (20584,-0.974593), (20585,-0.612235), (20586,-0.773359), (20587,-0.471845), (20588,-0.632499), (20589,-0.683073), (20590,-0.846520), (20591,-0.870613), (20592,-1.006659), (20593,-0.642898), (20594,-0.824459), (20595,-0.572645), (20596,-0.715190), (20597,-0.666360), (20598,-0.803332), (20599,-0.665787), (20600,-1.082380), (20601,-0.739527), (20602,-0.891358), (20603,-0.611673), (20604,-0.787662), (20605,-0.871216), (20606,-0.983567), (20607,-1.014167), (20608,-1.061021), (20609,-1.219822), (20610,-0.679557), (20611,-0.798877), (20612,-0.849915), (20613,-0.994313), (20614,-0.633345), (20615,-0.778677), (20616,-1.066142), (20617,-0.728862), (20618,-0.910887), (20619,-0.905719), (20620,-1.058947), (20621,-1.128563), (20622,-1.270181), (20623,-1.013257), (20624,-1.167412), (20625,-0.827345), (20626,-0.948056), (20627,-0.781713), (20628,-0.950732), (20629,-0.895866), (20630,-1.084854), (20631,-0.814461), (20632,-0.964439), (20633,-1.014079), (20634,-0.799428), (20635,-0.775682), (20636,-0.935879), (20637,-0.995739), (20638,-1.140607), (20639,-0.832124), (20640,-0.993248), (20641,-1.060077), (20642,-0.815231), (20643,-0.684649), (20644,-0.856925), (20645,-0.894023), (20646,-0.925092), (20647,-0.650053), (20648,-1.082438), (20649,-0.721470), (20650,-0.890953), (20651,-0.869530), (20652,-1.025081), (20653,-1.105379), (20654,-1.261393), (20655,-0.989140), (20656,-1.148874), (20657,-0.833891), (20658,-0.959712), (20659,-0.842598), (20660,-1.003258), (20661,-0.949782), (20662,-1.083035), (20663,-0.820074), (20664,-0.985381), (20665,-1.069862), (20666,-0.826876), (20667,-0.801734), (20668,-0.962394), (20669,-1.011108), (20670,-1.187560), (20671,-0.909271), (20672,-1.072718), (20673,-1.146516), (20674,-0.929072), (20675,-0.740431), (20676,-0.920596), (20677,-0.944696), (20678,-1.015708), (20679,-0.746705), (20680,-1.073193), (20681,-0.728943), (20682,-0.887281), (20683,-0.843560), (20684,-0.980526), (20685,-1.075226), (20686,-1.233100), (20687,-0.968743), (20688,-1.167956), (20689,-0.812561), (20690,-0.971362), (20691,-0.811055), (20692,-0.926656), (20693,-0.910343), (20694,-1.045456), (20695,-0.808043), (20696,-0.951978), (20697,-1.006728), (20698,-0.798583), (20699,-0.792019), (20700,-0.946643), (20701,-0.998143), (20702,-1.181095), (20703,-0.864716), (20704,-1.016091), (20705,-1.087096), (20706,-0.845037), (20707,-0.657329), (20708,-0.810557), (20709,-0.885282), (20710,-0.933070), (20711,-0.661743), (20712,-0.842378), (20713,-0.898989), (20714,-0.653680), (20715,-0.618318), (20716,-0.804063), (20717,-0.865319), (20718,-1.051521), (20719,-0.732362), (20720,-0.905095), (20721,-0.968674), (20722,-0.734511), (20723,-0.569095), (20724,-0.706994), (20725,-0.779859), (20726,-0.860627), (20727,-0.592093), (20728,-0.782014), (20729,-0.839551), (20730,-0.628619), (20731,-0.587685), (20732,-0.765527), (20733,-0.801705), (20734,-0.989767), (20735,-0.724946), (20736,-0.892106), (20737,-0.935248), (20738,-0.686689), (20739,-0.525449), (20740,-0.663348), (20741,-0.724141), (20742,-0.803049), (20743,-0.515468), (20744,-0.804329), (20745,-0.892993), (20746,-0.661616), (20747,-0.626725), (20748,-0.791098), (20749,-0.852354), (20750,-1.025551), (20751,-0.762590), (20752,-0.914891), (20753,-0.964995), (20754,-0.726192), (20755,-0.554270), (20756,-0.723753), (20757,-0.785942), (20758,-0.824901), (20759,-0.557757), (20760,-0.929762), (20761,-1.086239), (20762,-0.678822), (20763,-0.803716), (20764,-0.875654), (20765,-1.042814), (20766,-0.767311), (20767,-0.942837), (20768,-1.004093), (20769,-1.137346), (20770,-0.574320), (20771,-0.747523), (20772,-0.781835), (20773,-0.946678), (20774,-0.601502), (20775,-0.740791), (20776,-0.827595), (20777,-0.985932), (20778,-0.578515), (20779,-0.718267), (20780,-0.802285), (20781,-0.976877), (20782,-0.713453), (20783,-0.884333), (20784,-0.920505), (20785,-1.065367), (20786,-0.545077), (20787,-0.679726), (20788,-0.757701), (20789,-0.890954), (20790,-0.511870), (20791,-0.672994), (20792,-0.880567), (20793,-1.023112), (20794,-0.653315), (20795,-0.789818), (20796,-0.836679), (20797,-1.009875), (20798,-0.745061), (20799,-0.901538), (20800,-0.946070), (20801,-1.081182), (20802,-0.546953), (20803,-0.696468), (20804,-0.727067), (20805,-0.872399), (20806,-0.529076), (20807,-0.700419), (20808,-0.815557), (20809,-0.973431), (20810,-0.579945), (20811,-0.754538), (20812,-0.810221), (20813,-0.925823), (20814,-0.657753), (20815,-0.815163), (20816,-0.932155), (20817,-1.023141), (20818,-0.460115), (20819,-0.604984), (20820,-0.695037), (20821,-0.831540), (20822,-0.464535), (20823,-0.659103), (20824,-0.900583), (20825,-1.051951), (20826,-0.640350), (20827,-0.772677), (20828,-0.850652), (20829,-0.979728), (20830,-0.749741), (20831,-0.897396), (20832,-0.936355), (20833,-1.103521), (20834,-0.551177), (20835,-0.730879), (20836,-0.786563), (20837,-0.943503), (20838,-0.573712), (20839,-0.720434), (20840,-0.984675), (20841,-0.648791), (20842,-0.806659), (20843,-0.775480), (20844,-0.930568), (20845,-0.994610), (20846,-1.142729), (20847,-0.902060), (20848,-1.055751), (20849,-0.720330), (20850,-0.851260), (20851,-0.740652), (20852,-0.888307), (20853,-0.832977), (20854,-0.999674), (20855,-0.732994), (20856,-0.928494), (20857,-1.051528), (20858,-0.665939), (20859,-0.817307), (20860,-0.867881), (20861,-1.037827), (20862,-0.775330), (20863,-0.915552), (20864,-1.068316), (20865,-1.104952), (20866,-0.884264), (20867,-0.748108), (20868,-0.885074), (20869,-0.950977), (20870,-1.031745), (20871,-0.770637), (20872,-1.005154), (20873,-1.071983), (20874,-0.815059), (20875,-0.803392), (20876,-0.949187), (20877,-1.020199), (20878,-1.192932), (20879,-0.904423), (20880,-1.058115), (20881,-1.130523), (20882,-0.907505), (20883,-0.733260), (20884,-0.870696), (20885,-0.943104), (20886,-1.036871), (20887,-0.736291), (20888,-0.890908), (20889,-1.040417), (20890,-0.692454), (20891,-0.825243), (20892,-0.821936), (20893,-0.946366), (20894,-1.035956), (20895,-1.192434), (20896,-0.938759), (20897,-1.055757), (20898,-0.714294), (20899,-0.876351), (20900,-0.749951), (20901,-0.897136), (20902,-0.862244), (20903,-1.024758), (20904,-1.017267), (20905,-0.792396), (20906,-0.827178), (20907,-0.967401), (20908,-0.938082), (20909,-1.129393), (20910,-1.163248), (20911,-1.335518), (20912,-1.066051), (20913,-0.851863), (20914,-0.913119), (20915,-1.060311), (20916,-0.914863), (20917,-0.958937), (20918,-1.000219), (20919,-1.178994), (20920,-0.909064), (20921,-1.073901), (20922,-0.724548), (20923,-0.879166), (20924,-0.874462), (20925,-1.008184), (20926,-1.104738), (20927,-1.237064), (20928,-0.958311), (20929,-1.096674), (20930,-0.772399), (20931,-0.923767), (20932,-0.795044), (20933,-0.942236), (20934,-0.892942), (20935,-1.056852), (20936,-0.811074), (20937,-0.979167), (20938,-0.633527), (20939,-0.777462), (20940,-0.771368), (20941,-0.912054), (20942,-1.019759), (20943,-1.165554), (20944,-0.884942), (20945,-1.066034), (20946,-0.694383), (20947,-0.833673), (20948,-0.694267), (20949,-0.868866), (20950,-0.850693), (20951,-0.998342), (20952,-0.882631), (20953,-1.015414), (20954,-0.666061), (20955,-0.816966), (20956,-0.806225), (20957,-0.940405), (20958,-1.029995), (20959,-1.199015), (20960,-0.900751), (20961,-1.030754), (20962,-0.680932), (20963,-0.842519), (20964,-0.730057), (20965,-0.904650), (20966,-0.872081), (20967,-1.041564), (20968,-0.768848), (20969,-0.890949), (20970,-0.538346), (20971,-0.678562), (20972,-0.698479), (20973,-0.838238), (20974,-0.913890), (20975,-1.078733), (20976,-0.807413), (20977,-0.927191), (20978,-0.600599), (20979,-0.737102), (20980,-0.625104), (20981,-0.821525), (20982,-0.797779), (20983,-0.960293), (20984,-0.816711), (20985,-0.897479), (20986,-0.580636), (20987,-0.765911), (20988,-0.740306), (20989,-0.896783), (20990,-0.954790), (20991,-1.109871), (20992,-0.851093), (20993,-0.991315), (20994,-0.666577), (20995,-0.823518), (20996,-0.679930), (20997,-0.835481), (20998,-0.797802), (20999,-0.942201), (21000,-0.834843), (21001,-0.997827), (21002,-0.644754), (21003,-0.807268), (21004,-0.797461), (21005,-1.008747), (21006,-1.063034), (21007,-1.208829), (21008,-0.940295), (21009,-1.074481), (21010,-0.717226), (21011,-0.875094), (21012,-0.726402), (21013,-0.872661), (21014,-0.834983), (21015,-0.994710), (21016,-0.960745), (21017,-1.013642), (21018,-0.747895), (21019,-0.763166), (21020,-0.904314), (21021,-0.970217), (21022,-1.147133), (21023,-0.871630), (21024,-1.037393), (21025,-1.062420), (21026,-0.844981), (21027,-0.680029), (21028,-0.841152), (21029,-0.884757), (21030,-0.967848), (21031,-0.691882), (21032,-0.860431), (21033,-0.919365), (21034,-0.727011), (21035,-0.706051), (21036,-0.810507), (21037,-0.866654), (21038,-1.038460), (21039,-0.779676), (21040,-0.964494), (21041,-1.000666), (21042,-0.761856), (21043,-0.591794), (21044,-0.724120), (21045,-0.799778), (21046,-0.902837), (21047,-0.591105), (21048,-0.955676), (21049,-1.040620), (21050,-0.775800), (21051,-0.739512), (21052,-0.882521), (21053,-0.916839), (21054,-1.101188), (21055,-0.830331), (21056,-1.038831), (21057,-1.073143), (21058,-0.812975), (21059,-0.658704), (21060,-0.810072), (21061,-0.896413), (21062,-0.928402), (21063,-0.640827), (21064,-0.903208), (21065,-0.998371), (21066,-0.746557), (21067,-0.749755), (21068,-0.906232), (21069,-0.980957), (21070,-1.155550), (21071,-0.839641), (21072,-1.015160), (21073,-1.049015), (21074,-0.811132), (21075,-0.649899), (21076,-0.811949), (21077,-0.895967), (21078,-0.975802), (21079,-0.662679), (21080,-0.954321), (21081,-0.988639), (21082,-0.725215), (21083,-0.712152), (21084,-0.859800), (21085,-0.930812), (21086,-1.112374), (21087,-0.842444), (21088,-0.961765), (21089,-1.025344), (21090,-0.792108), (21091,-0.655959), (21092,-0.809650), (21093,-0.848145), (21094,-0.928906), (21095,-0.665019), (21096,-1.018445), (21097,-0.676055), (21098,-0.811161), (21099,-0.792995), (21100,-0.955972), (21101,-1.052995), (21102,-1.222014), (21103,-0.959054), (21104,-1.095557), (21105,-0.748990), (21106,-0.895712), (21107,-0.773958), (21108,-0.908138), (21109,-0.871387), (21110,-1.017182), (21111,-0.742612), (21112,-0.909309), (21113,-0.948267), (21114,-0.734542), (21115,-0.699187), (21116,-0.877493), (21117,-0.959187), (21118,-1.144462), (21119,-0.856887), (21120,-1.135060), (21121,-1.171702), (21122,-0.917100), (21123,-0.761440), (21124,-0.943465), (21125,-0.965235), (21126,-1.055289), (21127,-0.733343), (21128,-0.911649), (21129,-1.045829), (21130,-0.683934), (21131,-0.874318), (21132,-0.867297), (21133,-1.001940), (21134,-1.075739), (21135,-1.221534), (21136,-0.952074), (21137,-1.114587), (21138,-0.769874), (21139,-0.911487), (21140,-0.774874), (21141,-0.929955), (21142,-0.902496), (21143,-1.073833), (21144,-1.017576), (21145,-1.161975), (21146,-0.778246), (21147,-0.932863), (21148,-0.927702), (21149,-1.112977), (21150,-1.196995), (21151,-1.350686), (21152,-1.052885), (21153,-1.216795), (21154,-0.863723), (21155,-1.016951), (21156,-0.875686), (21157,-1.020554), (21158,-0.968474), (21159,-1.113799), (21160,-0.886142), (21161,-1.048662), (21162,-0.745289), (21163,-0.873896), (21164,-0.854796), (21165,-1.006627), (21166,-1.109223), (21167,-1.267560), (21168,-1.001813), (21169,-1.110445), (21170,-0.803822), (21171,-0.947758), (21172,-0.791634), (21173,-0.938819), (21174,-0.910433), (21175,-1.012096), (21176,-0.913103), (21177,-1.083050), (21178,-0.758312), (21179,-0.900857), (21180,-0.923097), (21181,-1.061459), (21182,-1.172414), (21183,-1.327502), (21184,-1.019946), (21185,-1.199648), (21186,-0.856331), (21187,-1.042076), (21188,-0.890128), (21189,-1.012229), (21190,-0.986166), (21191,-1.143571), (21192,-0.914054), (21193,-1.058452), (21194,-0.697021), (21195,-0.848389), (21196,-0.835325), (21197,-1.012704), (21198,-1.103228), (21199,-1.255059), (21200,-0.970734), (21201,-1.130461), (21202,-0.747195), (21203,-0.920397), (21204,-0.756371), (21205,-0.912849), (21206,-0.901645), (21207,-1.058122), (21208,-1.021371), (21209,-1.159270), (21210,-0.798765), (21211,-0.931091), (21212,-0.947289), (21213,-1.088901), (21214,-1.190570), (21215,-1.338225), (21216,-1.065509), (21217,-1.201548), (21218,-0.847086), (21219,-1.010063), (21220,-0.851616), (21221,-1.023885), (21222,-0.982024), (21223,-1.147794), (21224,-0.836988), (21225,-1.006935), (21226,-0.692415), (21227,-0.826601), (21228,-0.798209), (21229,-0.937499), (21230,-1.027089), (21231,-1.174744), (21232,-0.915496), (21233,-1.089162), (21234,-0.728657), (21235,-0.858197), (21236,-0.712749), (21237,-0.878982), (21238,-0.864529), (21239,-1.024256), (21240,-0.792416), (21241,-0.928456), (21242,-0.587462), (21243,-0.768554), (21244,-0.755960), (21245,-0.917547), (21246,-0.996455), (21247,-1.161755), (21248,-0.900191), (21249,-1.043200), (21250,-0.718455), (21251,-0.880975), (21252,-0.703944), (21253,-0.871573), (21254,-0.838998), (21255,-0.995476), (21256,-0.855144), (21257,-0.994897), (21258,-0.644147), (21259,-0.785296), (21260,-0.781062), (21261,-0.911992), (21262,-1.005765), (21263,-1.177571), (21264,-0.910891), (21265,-1.071088), (21266,-0.733807), (21267,-0.879139), (21268,-0.715576), (21269,-0.881346), (21270,-0.854814), (21271,-0.994103), (21272,-0.851911), (21273,-0.917351), (21274,-1.051530), (21275,-0.642716), (21276,-0.753678), (21277,-0.833976), (21278,-0.964443), (21279,-0.729816), (21280,-0.896976), (21281,-0.951269), (21282,-1.087309), (21283,-0.565622), (21284,-0.725819), (21285,-0.807977), (21286,-0.935194), (21287,-0.563536), (21288,-0.949010), (21289,-1.013985), (21290,-0.787255), (21291,-0.761186), (21292,-0.910694), (21293,-0.964518), (21294,-1.131684), (21295,-0.845499), (21296,-0.992684), (21297,-1.053940), (21298,-0.808168), (21299,-0.691987), (21300,-0.802016), (21301,-0.879991), (21302,-0.953789), (21303,-0.665751), (21304,-0.931845), (21305,-0.968950), (21306,-0.758938), (21307,-0.767709), (21308,-0.985501), (21309,-1.035142), (21310,-1.202308), (21311,-0.891038), (21312,-1.050302), (21313,-1.111095), (21314,-0.880182), (21315,-0.730094), (21316,-0.867530), (21317,-0.906489), (21318,-0.961245), (21319,-0.692242), (21320,-0.942551), (21321,-0.973150), (21322,-0.725055), (21323,-0.730569), (21324,-0.905162), (21325,-0.950626), (21326,-1.104317), (21327,-0.806987), (21328,-0.953708), (21329,-1.005209), (21330,-0.781728), (21331,-0.636287), (21332,-0.779295), (21333,-0.859130), (21334,-0.943147), (21335,-0.662072), (21336,-0.764204), (21337,-0.800840), (21338,-0.933629), (21339,-0.542004), (21340,-0.714743), (21341,-0.796437), (21342,-0.928757), (21343,-0.660224), (21344,-0.823207), (21345,-0.863562), (21346,-1.032576), (21347,-0.477915), (21348,-0.615351), (21349,-0.668241), (21350,-0.833085), (21351,-0.519492), (21352,-0.777697), (21353,-0.912803), (21354,-0.570883), (21355,-0.732470), (21356,-0.719870), (21357,-0.869848), (21358,-0.950609), (21359,-1.099191), (21360,-0.826474), (21361,-0.998750), (21362,-0.659610), (21363,-0.785430), (21364,-0.636269), (21365,-0.813648), (21366,-0.771324), (21367,-0.937094), (21368,-0.935176), (21369,-0.972745), (21370,-0.706534), (21371,-0.703690), (21372,-0.848088), (21373,-0.901449), (21374,-1.113204), (21375,-0.822836), (21376,-1.095906), (21377,-1.236592), (21378,-0.926249), (21379,-1.071581), (21380,-0.976765), (21381,-1.123957), (21382,-1.038433), (21383,-1.182832), (21384,-1.001624), (21385,-1.175283), (21386,-0.837539), (21387,-0.964756), (21388,-0.973990), (21389,-1.158802), (21390,-1.215412), (21391,-1.370030), (21392,-1.114965), (21393,-1.223140), (21394,-0.893756), (21395,-1.053020), (21396,-0.902469), (21397,-1.046404), (21398,-1.018939), (21399,-1.167057), (21400,-0.871116), (21401,-1.040136), (21402,-1.061912), (21403,-0.812421), (21404,-0.799827), (21405,-0.949798), (21406,-1.015701), (21407,-1.177288), (21408,-0.926406), (21409,-1.077774), (21410,-1.098618), (21411,-0.872814), (21412,-0.723196), (21413,-0.841120), (21414,-0.883328), (21415,-0.978028), (21416,-0.876713), (21417,-1.063847), (21418,-0.717281), (21419,-0.843101), (21420,-0.840720), (21421,-0.986052), (21422,-1.059850), (21423,-1.211218), (21424,-0.949648), (21425,-1.098229), (21426,-0.736798), (21427,-0.912780), (21428,-0.764552), (21429,-0.928463), (21430,-0.888925), (21431,-1.031933), (21432,-1.021656), (21433,-1.167915), (21434,-0.840853), (21435,-0.988039), (21436,-0.961043), (21437,-1.130063), (21438,-1.226159), (21439,-1.374740), (21440,-1.108524), (21441,-1.223198), (21442,-0.887314), (21443,-1.052151), (21444,-0.872803), (21445,-1.022774), (21446,-1.006461), (21447,-1.185700), (21448,-0.926452), (21449,-1.092686), (21450,-0.752619), (21451,-0.915602), (21452,-0.894643), (21453,-1.033469), (21454,-1.113303), (21455,-1.303694), (21456,-1.010540), (21457,-1.170267), (21458,-0.853425), (21459,-0.969489), (21460,-0.838450), (21461,-0.976812), (21462,-0.955853), (21463,-1.159243), (21464,-0.870271), (21465,-1.013743), (21466,-1.038306), (21467,-0.829227), (21468,-0.802695), (21469,-0.966605), (21470,-1.007886), (21471,-1.194558), (21472,-0.895361), (21473,-1.037443), (21474,-1.071292), (21475,-0.861749), (21476,-0.732100), (21477,-0.920161), (21478,-0.950297), (21479,-1.011553), (21480,-1.068633), (21481,-0.787088), (21482,-0.917091), (21483,-0.567268), (21484,-0.713064), (21485,-0.716262), (21486,-0.885745), (21487,-0.956757), (21488,-1.112765), (21489,-0.817757), (21490,-0.977021), (21491,-0.645313), (21492,-0.839880), (21493,-0.657276), (21494,-0.816077), (21495,-0.798837), (21496,-0.708667), (21497,-0.839597), (21498,-0.902249), (21499,-0.664836), (21500,-0.638304), (21501,-0.797568), (21502,-0.825844), (21503,-1.025057), (21504,-0.671052), (21505,-0.822883), (21506,-0.844197), (21507,-0.625362), (21508,-0.487816), (21509,-0.636398), (21510,-0.723202), (21511,-0.771916), (21512,-0.946045), (21513,-0.703059), (21514,-0.870683), (21515,-0.519470), (21516,-0.675015), (21517,-0.652202), (21518,-0.835154), (21519,-0.912665), (21520,-1.035236), (21521,-0.794110), (21522,-0.947337), (21523,-0.579400), (21524,-0.758169), (21525,-0.584857), (21526,-0.735761), (21527,-0.694364), (21528,-0.820184), (21529,-0.900025), (21530,-1.043960), (21531,-0.633757), (21532,-0.764223), (21533,-0.818510), (21534,-0.971268), (21535,-0.732002), (21536,-0.879650), (21537,-0.923725), (21538,-1.054655), (21539,-0.520889), (21540,-0.652752), (21541,-0.726551), (21542,-0.929940), (21543,-0.567576), (21544,-0.680860), (21545,-0.825259), (21546,-0.874437), (21547,-0.633774), (21548,-0.590986), (21549,-0.756286), (21550,-0.816616), (21551,-0.988885), (21552,-0.731498), (21553,-0.893085), (21554,-0.922757), (21555,-0.668156), (21556,-0.529214), (21557,-0.675472), (21558,-0.750667), (21559,-0.836544), (21560,-0.740332), (21561,-0.800662), (21562,-0.932055), (21563,-0.551582), (21564,-0.727564), (21565,-0.759560), (21566,-0.917427), (21567,-0.662832), (21568,-0.822096), (21569,-0.857805), (21570,-1.025898), (21571,-0.479127), (21572,-0.640251), (21573,-0.708940), (21574,-0.856125), (21575,-0.484011), (21576,-0.634452), (21577,-0.790930), (21578,-0.850789), (21579,-0.586902), (21580,-0.590094), (21581,-0.759577), (21582,-0.797145), (21583,-0.975921), (21584,-0.692059), (21585,-0.868974), (21586,-0.943699), (21587,-0.690495), (21588,-0.550626), (21589,-0.696421), (21590,-0.728410), (21591,-0.798959), (21592,-0.819802), (21593,-0.854121), (21594,-1.016171), (21595,-0.606894), (21596,-0.773591), (21597,-0.815805), (21598,-0.950448), (21599,-0.646612), (21600,-0.855117), (21601,-0.895472), (21602,-1.041731), (21603,-0.513544), (21604,-0.658870), (21605,-0.702474), (21606,-0.870104), (21607,-0.474296), (21608,-0.674899), (21609,-0.812799), (21610,-0.507108), (21611,-0.652434), (21612,-0.637047), (21613,-0.754978), (21614,-0.848281), (21615,-1.019624), (21616,-0.734829), (21617,-0.892703), (21618,-0.557746), (21619,-0.702608), (21620,-0.551130), (21621,-0.706681), (21622,-0.685252), (21623,-0.823614), (21624,-0.791046), (21625,-0.962852), (21626,-0.643686), (21627,-0.788555), (21628,-0.774095), (21629,-0.968662), (21630,-1.041534), (21631,-1.198011), (21632,-0.915539), (21633,-1.078060), (21634,-1.117481), (21635,-0.900506), (21636,-0.745309), (21637,-0.927334), (21638,-0.948178), (21639,-0.992715), (21640,-0.955494), (21641,-1.129624), (21642,-0.787234), (21643,-0.948821), (21644,-0.937154), (21645,-1.078303), (21646,-1.160930), (21647,-1.323444), (21648,-1.050727), (21649,-1.213711), (21650,-0.817903), (21651,-0.957192), (21652,-0.840548), (21653,-0.957082), (21654,-0.937513), (21655,-1.123721), (21656,-0.769722), (21657,-0.939668), (21658,-0.986059), (21659,-0.766761), (21660,-0.755094), (21661,-0.887884), (21662,-0.937061), (21663,-1.113050), (21664,-0.844047), (21665,-1.018176), (21666,-1.092901), (21667,-0.859208), (21668,-0.705864), (21669,-0.852592), (21670,-0.906416), (21671,-0.989500), (21672,-1.303910), (21673,-1.009828), (21674,-0.757087), (21675,-0.864329), (21676,-1.022197), (21677,-1.023998), (21678,-1.211596), (21679,-1.230586), (21680,-1.375918), (21681,-1.100879), (21682,-0.847674), (21683,-0.900564), (21684,-1.034750), (21685,-0.892559), (21686,-0.984002), (21687,-1.002066), (21688,-1.192450), (21689,-0.916948), (21690,-1.083644), (21691,-0.760302), (21692,-0.900982), (21693,-0.866553), (21694,-1.023964), (21695,-1.110304), (21696,-1.259349), (21697,-0.974091), (21698,-1.145897), (21699,-0.801647), (21700,-0.946052), (21701,-0.758338), (21702,-0.944077), (21703,-0.908258), (21704,-1.200363), (21705,-0.946695), (21706,-0.682345), (21707,-0.748710), (21708,-0.920516), (21709,-0.903733), (21710,-1.065784), (21711,-1.135406), (21712,-1.311858), (21713,-1.017307), (21714,-0.781754), (21715,-0.828145), (21716,-1.024109), (21717,-0.874484), (21718,-0.961752), (21719,-1.022075), (21720,-1.189705), (21721,-0.927671), (21722,-1.096227), (21723,-0.751514), (21724,-0.873621), (21725,-0.875886), (21726,-1.037473), (21727,-1.136356), (21728,-1.274719), (21729,-0.955090), (21730,-1.117140), (21731,-0.777073), (21732,-0.929368), (21733,-0.799255), (21734,-0.957592), (21735,-0.900866), (21736,-1.042942), (21737,-0.789737), (21738,-0.955970), (21739,-0.585246), (21740,-0.720359), (21741,-0.702649), (21742,-0.863773), (21743,-0.938962), (21744,-1.107054), (21745,-0.818083), (21746,-0.967128), (21747,-0.630311), (21748,-0.788648), (21749,-0.651566), (21750,-0.808970), (21751,-0.796840), (21752,-0.999766), (21753,-0.709862), (21754,-0.867736), (21755,-0.507694), (21756,-0.659062), (21757,-0.643212), (21758,-0.827097), (21759,-0.887426), (21760,-1.055513), (21761,-0.799058), (21762,-0.932311), (21763,-0.583416), (21764,-0.718992), (21765,-0.579586), (21766,-0.750929), (21767,-0.707678), (21768,-0.993747), (21769,-0.702916), (21770,-0.895623), (21771,-0.553234), (21772,-0.720400), (21773,-0.709196), (21774,-0.872636), (21775,-0.935752), (21776,-1.079688), (21777,-0.831129), (21778,-0.960199), (21779,-0.597371), (21780,-0.763141), (21781,-0.651607), (21782,-0.804834), (21783,-0.769473), (21784,-0.786140), (21785,-0.941221), (21786,-1.008520), (21787,-0.789685), (21788,-0.787304), (21789,-0.944245), (21790,-0.986460), (21791,-1.149443), (21792,-0.834454), (21793,-1.014626), (21794,-1.068913), (21795,-0.825927), (21796,-0.696271), (21797,-0.854608), (21798,-0.897750), (21799,-0.954360), (21800,-0.708588), (21801,-0.852986), (21802,-0.920285), (21803,-0.652215), (21804,-0.629396), (21805,-0.804921), (21806,-0.848989), (21807,-1.040770), (21808,-0.790352), (21809,-0.911989), (21810,-0.975105), (21811,-0.732119), (21812,-0.575989), (21813,-0.735723), (21814,-0.813698), (21815,-0.878674), (21816,-0.669125), (21817,-0.829322), (21818,-0.912870), (21819,-0.680566), (21820,-0.632669), (21821,-0.804012), (21822,-0.865732), (21823,-1.019886), (21824,-0.776900), (21825,-0.933378), (21826,-0.978842), (21827,-0.798561), (21828,-0.639180), (21829,-0.793805), (21830,-0.850415), (21831,-0.936755), (21832,-0.717921), (21833,-0.862783), (21834,-0.903601), (21835,-0.690346), (21836,-0.681459), (21837,-0.838869), (21838,-0.886187), (21839,-1.040348), (21840,-0.749053), (21841,-0.881373), (21842,-0.950062), (21843,-0.746556), (21844,-0.583463), (21845,-0.757128), (21846,-0.818385), (21847,-0.888927), (21848,-0.790868), (21849,-0.945485), (21850,-1.004419), (21851,-0.798590), (21852,-0.785996), (21853,-0.955009), (21854,-1.002333), (21855,-1.176462), (21856,-0.898636), (21857,-1.036536), (21858,-1.073171), (21859,-0.845514), (21860,-0.674525), (21861,-0.823106), (21862,-0.849992), (21863,-0.934936), (21864,-0.873564), (21865,-0.995671), (21866,-0.675579), (21867,-0.824161), (21868,-0.835712), (21869,-0.999159), (21870,-1.076670), (21871,-1.252659), (21872,-0.967401), (21873,-1.104836), (21874,-0.784744), (21875,-0.930539), (21876,-0.806463), (21877,-0.957831), (21878,-0.914573), (21879,-1.039930), (21880,-0.797408), (21881,-0.937630), (21882,-0.983558), (21883,-0.717348), (21884,-0.666658), (21885,-0.801770), (21886,-0.891824), (21887,-1.039016), (21888,-0.973460), (21889,-1.143413), (21890,-0.785225), (21891,-0.948672), (21892,-0.781865), (21893,-0.936947), (21894,-0.919707), (21895,-1.085933), (21896,-0.889397), (21897,-1.041698), (21898,-0.717886), (21899,-0.849279), (21900,-0.821820), (21901,-0.985267), (21902,-1.095296), (21903,-1.255950), (21904,-0.974411), (21905,-1.115560), (21906,-0.768993), (21907,-0.952872), (21908,-0.810680), (21909,-0.965304), (21910,-0.916474), (21911,-1.070628), (21912,-1.092405), (21913,-0.810860), (21914,-0.985458), (21915,-0.630526), (21916,-0.776322), (21917,-0.757215), (21918,-0.920199), (21919,-1.010253), (21920,-1.156981), (21921,-0.902379), (21922,-1.053284), (21923,-0.728076), (21924,-0.865512), (21925,-0.706602), (21926,-0.859823), (21927,-0.849083), (21928,-1.189503), (21929,-0.902391), (21930,-0.668228), (21931,-0.742026), (21932,-0.897108), (21933,-0.866862), (21934,-1.051204), (21935,-1.113393), (21936,-1.262438), (21937,-0.990655), (21938,-0.755095), (21939,-0.813102), (21940,-0.970043), (21941,-0.823675), (21942,-0.897936), (21943,-0.948041), (21944,-1.352562), (21945,-1.045475), (21946,-0.793660), (21947,-0.850270), (21948,-1.044838), (21949,-1.022019), (21950,-1.226805), (21951,-1.269019), (21952,-1.414351), (21953,-1.149068), (21954,-0.911185), (21955,-0.956186), (21956,-1.122419), (21957,-0.978831), (21958,-1.025228), (21959,-1.075333), (21960,-1.298697), (21961,-0.991611), (21962,-0.756984), (21963,-0.798735), (21964,-0.961712), (21965,-0.952368), (21966,-1.124638), (21967,-1.192863), (21968,-1.361883), (21969,-1.104495), (21970,-0.845248), (21971,-0.898608), (21972,-1.070878), (21973,-0.938905), (21974,-0.975547), (21975,-1.017292), (21976,-1.184921), (21977,-0.886194), (21978,-1.056140), (21979,-0.692849), (21980,-0.844217), (21981,-0.800960), (21982,-0.965339), (21983,-1.063289), (21984,-1.214194), (21985,-0.960983), (21986,-1.085876), (21987,-0.759748), (21988,-0.915762), (21989,-0.775424), (21990,-0.919359), (21991,-0.894687), (21992,-1.064633), (21993,-0.759406), (21994,-0.922853), (21995,-0.588822), (21996,-0.730898), (21997,-0.752674), (21998,-0.892897), (21999,-0.945324), (22000,-1.091582), (22001,-0.847670), (22002,-1.009720), (22003,-0.670580), (22004,-0.791297), (22005,-0.607760), (22006,-0.758664), (22007,-0.754893), (22008,-0.975935), (22009,-0.666062), (22010,-0.824399), (22011,-0.449492), (22012,-0.656138), (22013,-0.613344), (22014,-0.779114), (22015,-0.876601), (22016,-1.087423), (22017,-0.814243), (22018,-0.963295), (22019,-0.637623), (22020,-0.770876), (22021,-0.623575), (22022,-0.755901), (22023,-0.721936), (22024,-1.003829), (22025,-0.707425), (22026,-0.875048), (22027,-0.525689), (22028,-0.697965), (22029,-0.692334), (22030,-0.835336), (22031,-0.903098), (22032,-1.048894), (22033,-0.770604), (22034,-0.917790), (22035,-0.581906), (22036,-0.723054), (22037,-0.601764), (22038,-0.763351), (22039,-0.709412), (22040,-0.746980), (22041,-0.899744), (22042,-0.939166), (22043,-0.719868), (22044,-0.696122), (22045,-0.885117), (22046,-0.898064), (22047,-1.066157), (22048,-0.764180), (22049,-0.916938), (22050,-0.980517), (22051,-0.715234), (22052,-0.604163), (22053,-0.743458), (22054,-0.825152), (22055,-0.896628), (22056,-0.605797), (22057,-0.774353), (22058,-0.865797), (22059,-0.618165), (22060,-0.618107), (22061,-0.769011), (22062,-0.810762), (22063,-0.985818), (22064,-0.718675), (22065,-0.845892), (22066,-0.871845), (22067,-0.646047), (22068,-0.500606), (22069,-0.694240), (22070,-0.736454), (22071,-0.777736), (22072,-0.629502), (22073,-0.805027), (22074,-0.847705), (22075,-0.605183), (22076,-0.588400), (22077,-0.752310), (22078,-0.823322), (22079,-1.009993), (22080,-0.700120), (22081,-0.860311), (22082,-0.901592), (22083,-0.692513), (22084,-0.534066), (22085,-0.662210), (22086,-0.713710), (22087,-0.813983), (22088,-0.615123), (22089,-0.778107), (22090,-0.808706), (22091,-0.568043), (22092,-0.591210), (22093,-0.765339), (22094,-0.763891), (22095,-0.950092), (22096,-0.674126), (22097,-0.867297), (22098,-0.896970), (22099,-0.637259), (22100,-0.476489), (22101,-0.644582), (22102,-0.697472), (22103,-0.786136), (22104,-0.708972), (22105,-0.881248), (22106,-0.929029), (22107,-0.704158), (22108,-0.700850), (22109,-0.860114), (22110,-0.921370), (22111,-1.115474), (22112,-0.832075), (22113,-0.972298), (22114,-0.992214), (22115,-0.742723), (22116,-0.597745), (22117,-0.776983), (22118,-0.827551), (22119,-0.886021), (22120,-0.727574), (22121,-0.891947), (22122,-0.536088), (22123,-0.692566), (22124,-0.713879), (22125,-0.840626), (22126,-0.920461), (22127,-1.057897), (22128,-0.782857), (22129,-0.932835), (22130,-0.602987), (22131,-0.753422), (22132,-0.588939), (22133,-0.713833), (22134,-0.703556), (22135,-0.856783), (22136,-0.805167), (22137,-0.952352), (22138,-0.632260), (22139,-0.801743), (22140,-0.809581), (22141,-0.945157), (22142,-1.030571), (22143,-1.175433), (22144,-0.920832), (22145,-1.069883), (22146,-1.111628), (22147,-0.890007), (22148,-0.736669), (22149,-0.886641), (22150,-0.940464), (22151,-1.047243), (22152,-1.324953), (22153,-1.019726), (22154,-0.775807), (22155,-0.863074), (22156,-1.036740), (22157,-1.030183), (22158,-1.215458), (22159,-1.208900), (22160,-1.334720), (22161,-1.062467), (22162,-0.838060), (22163,-0.909072), (22164,-1.044185), (22165,-0.880158), (22166,-0.946524), (22167,-1.031005), (22168,-1.173087), (22169,-0.895725), (22170,-1.078213), (22171,-0.765554), (22172,-0.920635), (22173,-0.887603), (22174,-1.021319), (22175,-1.109513), (22176,-1.269247), (22177,-1.013255), (22178,-1.156258), (22179,-0.795290), (22180,-0.981034), (22181,-0.835123), (22182,-0.973949), (22183,-0.924192), (22184,-1.331963), (22185,-1.042528), (22186,-0.782354), (22187,-0.842677), (22188,-1.029348), (22189,-1.016285), (22190,-1.180195), (22191,-1.189893), (22192,-1.358449), (22193,-1.075050), (22194,-0.850180), (22195,-0.898894), (22196,-1.074413), (22197,-0.895528), (22198,-0.967930), (22199,-1.015717), (22200,-1.242338), (22201,-0.946861), (22202,-1.140965), (22203,-0.801824), (22204,-0.941583), (22205,-0.928050), (22206,-1.057127), (22207,-1.159259), (22208,-1.332925), (22209,-1.055562), (22210,-1.190675), (22211,-0.869187), (22212,-1.023805), (22213,-0.865358), (22214,-0.986995), (22215,-0.961396), (22216,-1.262793), (22217,-0.994260), (22218,-0.742445), (22219,-0.803238), (22220,-0.963898), (22221,-0.955481), (22222,-1.140756), (22223,-1.176001), (22224,-1.323186), (22225,-1.050007), (22226,-0.780547), (22227,-0.826938), (22228,-1.001067), (22229,-0.867698), (22230,-0.896444), (22231,-0.947011), (22232,-1.138792), (22233,-0.867472), (22234,-1.021163), (22235,-0.699211), (22236,-0.808776), (22237,-0.797573), (22238,-0.940581), (22239,-1.042244), (22240,-1.187576), (22241,-0.939481), (22242,-1.101994), (22243,-0.747995), (22244,-0.928161), (22245,-0.785042), (22246,-0.941520), (22247,-0.907555), (22248,-1.039875), (22249,-0.768555), (22250,-0.903668), (22251,-0.553382), (22252,-0.720078), (22253,-0.744172), (22254,-0.917837), (22255,-0.969808), (22256,-1.097481), (22257,-0.851246), (22258,-0.979853), (22259,-0.638396), (22260,-0.816701), (22261,-0.655931), (22262,-0.812872), (22263,-0.742677), (22264,-0.966505), (22265,-0.667315), (22266,-0.846553), (22267,-0.475366), (22268,-0.623021), (22269,-0.624816), (22270,-0.776191), (22271,-0.871354), (22272,-1.025972), (22273,-0.771370), (22274,-0.931567), (22275,-0.568739), (22276,-0.713138), (22277,-0.588598), (22278,-0.741826), (22279,-0.717616), (22280,-1.022264), (22281,-0.717037), (22282,-0.884197), (22283,-0.551563), (22284,-0.711290), (22285,-0.714952), (22286,-0.860283), (22287,-0.925716), (22288,-1.053396), (22289,-0.819233), (22290,-0.955742), (22291,-0.598024), (22292,-0.723381), (22293,-0.578866), (22294,-0.751135), (22295,-0.746901), (22296,-0.738947), (22297,-0.888918), (22298,-0.962253), (22299,-0.730413), (22300,-0.724319), (22301,-0.878010), (22302,-0.911859), (22303,-1.081812), (22304,-0.816058), (22305,-1.008303), (22306,-1.021720), (22307,-0.787557), (22308,-0.626323), (22309,-0.794410), (22310,-0.864958), (22311,-0.925751), (22312,-0.715276), (22313,-0.873150), (22314,-0.901889), (22315,-0.644502), (22316,-0.641657), (22317,-0.813000), (22318,-0.834313), (22319,-1.033057), (22320,-0.766383), (22321,-0.922391), (22322,-0.979007), (22323,-0.753667), (22324,-0.552484), (22325,-0.710821), (22326,-0.752103), (22327,-0.833797), (22328,-0.651662), (22329,-0.799311), (22330,-0.859640), (22331,-0.599930), (22332,-0.595232), (22333,-0.772611), (22334,-0.806460), (22335,-0.992204), (22336,-0.710196), (22337,-0.846705), (22338,-0.904242), (22339,-0.666365), (22340,-0.536246), (22341,-0.713162), (22342,-0.781850), (22343,-0.851936), (22344,-0.675837), (22345,-0.817449), (22346,-0.890784), (22347,-0.655688), (22348,-0.624979), (22349,-0.774488), (22350,-0.829244), (22351,-0.989435), (22352,-0.714396), (22353,-0.870410), (22354,-0.932129), (22355,-0.700759), (22356,-0.534873), (22357,-0.683924), (22358,-0.742858), (22359,-0.826405), (22360,-0.716267), (22361,-0.846734), (22362,-0.894051), (22363,-0.662211), (22364,-0.669592), (22365,-0.824210), (22366,-0.870138), (22367,-1.080034), (22368,-0.811964), (22369,-0.939174), (22370,-1.025051), (22371,-0.768127), (22372,-0.628258), (22373,-0.802387), (22374,-0.853888), (22375,-0.906322), (22376,-0.825907), (22377,-0.983775), (22378,-0.628386), (22379,-0.764425), (22380,-0.756471), (22381,-0.899010), (22382,-0.943548), (22383,-1.094916), (22384,-0.838461), (22385,-1.004688), (22386,-0.641867), (22387,-0.794161), (22388,-0.658006), (22389,-0.812630), (22390,-0.794920), (22391,-0.939319), (22392,-0.726990), (22393,-0.912265), (22394,-0.977704), (22395,-0.758870), (22396,-0.745806), (22397,-0.906930), (22398,-0.956107), (22399,-1.105152), (22400,-0.936486), (22401,-1.089251), (22402,-1.154683), (22403,-0.884760), (22404,-0.751391), (22405,-0.912978), (22406,-0.948687), (22407,-1.015985), (22408,-1.157598), (22409,-0.869090), (22410,-1.030677), (22411,-0.695719), (22412,-0.864276), (22413,-0.848426), (22414,-1.010476), (22415,-1.069873), (22416,-1.213345), (22417,-0.947134), (22418,-1.099429), (22419,-0.757972), (22420,-0.894938), (22421,-0.742991), (22422,-0.887396), (22423,-0.858540), (22424,-1.137177), (22425,-0.860747), (22426,-1.008866), (22427,-0.690627), (22428,-0.810411), (22429,-0.810823), (22430,-0.941283), (22431,-1.016478), (22432,-1.167382), (22433,-0.896063), (22434,-1.055790), (22435,-0.725942), (22436,-0.875450), (22437,-0.726759), (22438,-0.853969), (22439,-0.828370), (22440,-1.265865), (22441,-1.016837), (22442,-0.779887), (22443,-0.844400), (22444,-1.006450), (22445,-0.993387), (22446,-1.140572), (22447,-1.180927), (22448,-1.356452), (22449,-1.083272), (22450,-0.812879), (22451,-0.881568), (22452,-1.028753), (22453,-0.913506), (22454,-0.952927), (22455,-0.953339), (22456,-1.159515), (22457,-0.917920), (22458,-1.050709), (22459,-0.718075), (22460,-0.842036), (22461,-0.872641), (22462,-1.022613), (22463,-1.085729), (22464,-1.268681), (22465,-1.013153), (22466,-1.166844), (22467,-0.853251), (22468,-0.987901), (22469,-0.829447), (22470,-0.971066), (22471,-0.944064), (22472,-1.120980), (22473,-0.858489), (22474,-1.020076), (22475,-0.665144), (22476,-0.807219), (22477,-0.786730), (22478,-0.928342), (22479,-1.026291), (22480,-1.173483), (22481,-0.918418), (22482,-1.057708), (22483,-0.700922), (22484,-0.873192), (22485,-0.756547), (22486,-0.893050), (22487,-0.862335), (22488,-1.177208), (22489,-0.911924), (22490,-1.089303), (22491,-0.771998), (22492,-0.880166), (22493,-0.878718), (22494,-1.060743), (22495,-1.147547), (22496,-1.304025), (22497,-1.023876), (22498,-1.184536), (22499,-0.863048), (22500,-0.985155), (22501,-0.854109), (22502,-1.004087), (22503,-0.955720), (22504,-1.095942), (22505,-0.793965), (22506,-0.990386), (22507,-0.604333), (22508,-0.772890), (22509,-0.775618), (22510,-0.922346), (22511,-0.994285), (22512,-1.134038), (22513,-0.849249), (22514,-0.995507), (22515,-0.654507), (22516,-0.805882), (22517,-0.676696), (22518,-0.871257), (22519,-0.815927), (22520,-1.102466), (22521,-0.810701), (22522,-0.949997), (22523,-0.620612), (22524,-0.769657), (22525,-0.790037), (22526,-0.937692), (22527,-1.000345), (22528,-1.250647), (22529,-0.960279), (22530,-1.105611), (22531,-1.163154), (22532,-0.951752), (22533,-0.769611), (22534,-0.923765), (22535,-0.956688), (22536,-1.199564), (22537,-0.922671), (22538,-1.084258), (22539,-1.126930), (22540,-0.867225), (22541,-0.870417), (22542,-1.036187), (22543,-1.069109), (22544,-1.260890), (22545,-0.981204), (22546,-1.133036), (22547,-1.175250), (22548,-0.957342), (22549,-0.816084), (22550,-0.983244), (22551,-1.041713), (22552,-0.897199), (22553,-1.044384), (22554,-1.089848), (22555,-1.215668), (22556,-0.811501), (22557,-0.960552), (22558,-1.013912), (22559,-1.173640), (22560,-0.913466), (22561,-1.062511), (22562,-1.135382), (22563,-1.291396), (22564,-0.759491), (22565,-0.913645), (22566,-0.984194), (22567,-1.142061), (22568,-0.883747), (22569,-1.002604), (22570,-1.052709), (22571,-1.209186), (22572,-0.815707), (22573,-0.943851), (22574,-0.988845), (22575,-1.134641), (22576,-0.900014), (22577,-1.060674), (22578,-1.127504), (22579,-1.283518), (22580,-0.761368), (22581,-0.909023), (22582,-0.946121), (22583,-1.120250), (22584,-0.861936), (22585,-0.976611), (22586,-1.071774), (22587,-1.198058), (22588,-0.824547), (22589,-0.951301), (22590,-0.982363), (22591,-1.133731), (22592,-0.869844), (22593,-1.028181), (22594,-1.078755), (22595,-1.255671), (22596,-0.718192), (22597,-0.883492), (22598,-0.951718), (22599,-1.126774), (22600,-0.877751), (22601,-1.025400), (22602,-1.105704), (22603,-1.283083), (22604,-0.858478), (22605,-1.006596), (22606,-1.030226), (22607,-1.187173), (22608,-0.941858), (22609,-1.095549), (22610,-1.148446), (22611,-1.290528), (22612,-0.734001), (22613,-0.842639), (22614,-0.921084), (22615,-1.067343), (22616,-0.791840), (22617,-0.917197), (22618,-1.000745), (22619,-1.146540), (22620,-0.754451), (22621,-0.912788), (22622,-0.966612), (22623,-1.103584), (22624,-0.886140), (22625,-1.028222), (22626,-1.110380), (22627,-1.266394), (22628,-0.719623), (22629,-0.862168), (22630,-0.935040), (22631,-1.101736), (22632,-0.960471), (22633,-1.092328), (22634,-1.127110), (22635,-0.910598), (22636,-0.867347), (22637,-1.038684), (22638,-1.073002), (22639,-1.305190), (22640,-1.004609), (22641,-1.161087), (22642,-1.193546), (22643,-0.941731), (22644,-0.797216), (22645,-0.930932), (22646,-1.006590), (22647,-1.051122), (22648,-1.025053), (22649,-1.209864), (22650,-1.272054), (22651,-1.020702), (22652,-1.004389), (22653,-1.184561), (22654,-1.237451), (22655,-1.403684), (22656,-1.191356), (22657,-1.338078), (22658,-1.388188), (22659,-1.167494), (22660,-0.977926), (22661,-1.158092), (22662,-1.230963), (22663,-1.294073), (22664,-1.278693), (22665,-1.432847), (22666,-1.043545), (22667,-1.173078), (22668,-1.190209), (22669,-1.341113), (22670,-1.420485), (22671,-1.556987), (22672,-1.275448), (22673,-1.413811), (22674,-1.073744), (22675,-1.259019), (22676,-1.113578), (22677,-1.281664), (22678,-1.248632), (22679,-1.422761), (22680,-1.401802), (22681,-1.120726), (22682,-1.304142), (22683,-0.978940), (22684,-1.106620), (22685,-1.101916), (22686,-1.272795), (22687,-1.354490), (22688,-1.492389), (22689,-1.217349), (22690,-1.345956), (22691,-1.016572), (22692,-1.174446), (22693,-1.014602), (22694,-1.154361), (22695,-1.115287), (22696,-1.567647), (22697,-1.287035), (22698,-1.016642), (22699,-1.091830), (22700,-1.272929), (22701,-1.227818), (22702,-1.421452), (22703,-1.463667), (22704,-1.625717), (22705,-1.376225), (22706,-1.144385), (22707,-1.184277), (22708,-1.333785), (22709,-1.177198), (22710,-1.221266), (22711,-1.267193), (22712,-1.477553), (22713,-1.188118), (22714,-1.343199), (22715,-1.012888), (22716,-1.110844), (22717,-1.108926), (22718,-1.263544), (22719,-1.315977), (22720,-1.455736), (22721,-1.213677), (22722,-1.399879), (22723,-1.039374), (22724,-1.209327), (22725,-1.049946), (22726,-1.174370), (22727,-1.162240), (22728,-1.493831), (22729,-1.223438), (22730,-0.957228), (22731,-0.998509), (22732,-1.167066), (22733,-1.147496), (22734,-1.314663), (22735,-1.376846), (22736,-1.552834), (22737,-1.239242), (22738,-1.006012), (22739,-1.065408), (22740,-1.205161), (22741,-1.064366), (22742,-1.152096), (22743,-1.188738), (22744,-1.360081), (22745,-1.084578), (22746,-1.256847), (22747,-0.943718), (22748,-1.105305), (22749,-1.120582), (22750,-1.286346), (22751,-1.348998), (22752,-1.474819), (22753,-1.198853), (22754,-1.380414), (22755,-1.018513), (22756,-1.160125), (22757,-1.018403), (22758,-1.173485), (22759,-1.133483), (22760,-1.311326), (22761,-1.055334), (22762,-1.202983), (22763,-0.850374), (22764,-1.016144), (22765,-1.024451), (22766,-1.159558), (22767,-1.222674), (22768,-1.364756), (22769,-1.122227), (22770,-1.283351), (22771,-0.954899), (22772,-1.095122), (22773,-0.926912), (22774,-1.107548), (22775,-1.078229), (22776,-1.250035), (22777,-0.988464), (22778,-1.132400), (22779,-0.805808), (22780,-0.958103), (22781,-0.942253), (22782,-1.074579), (22783,-1.158597), (22784,-1.218456), (22785,-0.942027), (22786,-1.105004), (22787,-0.773303), (22788,-0.938140), (22789,-0.775973), (22790,-0.942670), (22791,-0.935186), (22792,-1.238906), (22793,-0.956434), (22794,-1.090151), (22795,-0.768669), (22796,-0.905635), (22797,-0.933447), (22798,-1.078779), (22799,-1.137249), (22800,-1.261210), (22801,-0.991749), (22802,-1.169592), (22803,-0.832311), (22804,-0.966497), (22805,-0.832665), (22806,-0.969631), (22807,-0.941709), (22808,-0.968588), (22809,-1.138071), (22810,-1.201651), (22811,-0.982816), (22812,-0.980441), (22813,-1.142955), (22814,-1.176804), (22815,-1.345824), (22816,-1.075900), (22817,-1.205434), (22818,-1.244862), (22819,-1.029740), (22820,-0.876866), (22821,-0.998510), (22822,-1.033755), (22823,-1.100585), (22824,-0.855739), (22825,-1.034978), (22826,-1.068363), (22827,-0.839310), (22828,-0.841575), (22829,-1.012454), (22830,-1.082996), (22831,-1.243657), (22832,-0.972800), (22833,-1.105127), (22834,-1.155700), (22835,-0.935933), (22836,-0.763084), (22837,-0.898197), (22838,-0.965959), (22839,-1.043007), (22840,-0.889670), (22841,-1.056366), (22842,-1.134804), (22843,-0.873240), (22844,-0.873182), (22845,-1.087724), (22846,-1.098349), (22847,-1.248790), (22848,-0.989542), (22849,-1.132551), (22850,-1.190088), (22851,-0.947102), (22852,-0.809093), (22853,-0.961388), (22854,-0.992920), (22855,-1.078791), (22856,-0.899906), (22857,-1.022940), (22858,-1.082806), (22859,-0.863038), (22860,-0.869023), (22861,-0.999026), (22862,-1.057496), (22863,-1.238588), (22864,-0.937074), (22865,-1.098661), (22866,-1.152022), (22867,-0.939693), (22868,-0.758015), (22869,-0.938187), (22870,-0.956244), (22871,-1.033292), (22872,-0.898996), (22873,-1.080558), (22874,-1.154357), (22875,-0.880244), (22876,-0.860217), (22877,-1.051065), (22878,-1.084920), (22879,-1.265086), (22880,-0.966359), (22881,-1.130269), (22882,-1.159941), (22883,-0.946679), (22884,-0.769648), (22885,-0.910333), (22886,-0.979022), (22887,-1.065363), (22888,-1.024429), (22889,-1.151645), (22890,-0.800433), (22891,-0.973166), (22892,-0.946633), (22893,-1.117513), (22894,-1.205707), (22895,-1.345929), (22896,-1.079249), (22897,-1.251988), (22898,-0.894269), (22899,-1.049820), (22900,-0.928993), (22901,-1.053417), (22902,-1.044073), (22903,-1.150852), (22904,-0.957565), (22905,-1.135871), (22906,-1.148824), (22907,-0.912338), (22908,-0.925749), (22909,-1.049253), (22910,-1.081705), (22911,-1.286955), (22912,-1.107606), (22913,-1.281736), (22914,-1.345315), (22915,-1.090250), (22916,-0.951308), (22917,-1.103603), (22918,-1.114697), (22919,-1.168057), (22920,-1.171249), (22921,-1.310081), (22922,-0.985807), (22923,-1.152503), (22924,-1.148262), (22925,-1.279662), (22926,-1.348351), (22927,-1.494609), (22928,-1.220960), (22929,-1.377437), (22930,-1.055955), (22931,-1.184562), (22932,-1.056303), (22933,-1.220676), (22934,-1.154664), (22935,-1.321360), (22936,-1.310620), (22937,-1.028618), (22938,-1.167907), (22939,-0.841309), (22940,-1.023334), (22941,-0.995412), (22942,-1.185333), (22943,-1.225218), (22944,-1.345002), (22945,-1.090401), (22946,-1.241305), (22947,-0.917964), (22948,-1.064685), (22949,-0.955474), (22950,-1.098946), (22951,-1.062658), (22952,-1.513622), (22953,-1.252521), (22954,-0.999779), (22955,-1.022946), (22956,-1.181283), (22957,-1.161720), (22958,-1.352105), (22959,-1.420794), (22960,-1.598173), (22961,-1.325456), (22962,-1.082007), (22963,-1.088918), (22964,-1.240750), (22965,-1.102271), (22966,-1.184429), (22967,-1.249405), (22968,-1.437003), (22969,-1.165219), (22970,-1.331453), (22971,-0.967228), (22972,-1.087939), (22973,-1.120398), (22974,-1.257834), (22975,-1.343705), (22976,-1.489036), (22977,-1.228399), (22978,-1.373731), (22979,-1.041096), (22980,-1.202214), (22981,-1.037267), (22982,-1.147296), (22983,-1.121227), (22984,-1.426807), (22985,-1.144798), (22986,-0.930147), (22987,-0.973288), (22988,-1.122333), (22989,-1.128317), (22990,-1.308946), (22991,-1.388317), (22992,-1.540618), (22993,-1.273012), (22994,-1.023983), (22995,-1.081990), (22996,-1.198518), (22997,-1.016383), (22998,-1.131984), (22999,-1.212752), (23000,-1.351578), (23001,-1.093727), (23002,-1.229303), (23003,-0.889236), (23004,-1.030848), (23005,-1.046119), (23006,-1.211889), (23007,-1.340032), (23008,-1.476072), (23009,-1.193600), (23010,-1.321280), (23011,-0.987255), (23012,-1.139550), (23013,-1.008504), (23014,-1.175670), (23015,-1.139846), (23016,-1.301896), (23017,-1.007815), (23018,-1.168939), (23019,-0.809360), (23020,-0.981167), (23021,-0.973213), (23022,-1.087424), (23023,-1.183983), (23024,-1.313517), (23025,-1.050556), (23026,-1.207497), (23027,-0.863717), (23028,-0.995111), (23029,-0.839913), (23030,-0.984318), (23031,-0.937811), (23032,-1.229453), (23033,-0.969749), (23034,-1.113684), (23035,-0.780580), (23036,-0.926375), (23037,-0.949548), (23038,-1.103703), (23039,-1.170995), (23040,-1.335369), (23041,-1.055689), (23042,-1.194052), (23043,-0.841443), (23044,-0.980269), (23045,-0.837150), (23046,-1.033108), (23047,-1.042805), (23048,-1.347923), (23049,-1.125375), (23050,-1.237257), (23051,-0.881861), (23052,-1.081538), (23053,-1.076371), (23054,-1.219843), (23055,-1.296897), (23056,-1.439900), (23057,-1.187621), (23058,-1.332490), (23059,-0.993350), (23060,-1.172588), (23061,-1.027147), (23062,-1.189197), (23063,-1.145946), (23064,-1.059953), (23065,-1.249411), (23066,-1.244713), (23067,-1.012873), (23068,-0.971939), (23069,-1.146531), (23070,-1.164125), (23071,-1.334071), (23072,-1.047886), (23073,-1.179749), (23074,-1.195483), (23075,-0.970612), (23076,-0.832603), (23077,-1.002086), (23078,-1.067519), (23079,-1.156183), (23080,-0.911800), (23081,-1.060845), (23082,-1.111419), (23083,-0.891194), (23084,-0.884167), (23085,-1.032285), (23086,-1.072177), (23087,-1.285786), (23088,-1.007497), (23089,-1.146792), (23090,-1.208975), (23091,-0.926503), (23092,-0.788958), (23093,-0.952404), (23094,-0.970461), (23095,-1.067484), (23096,-0.973138), (23097,-1.119397), (23098,-1.190872), (23099,-0.939057), (23100,-0.879545), (23101,-1.057857), (23102,-1.120966), (23103,-1.250043), (23104,-1.014483), (23105,-1.160278), (23106,-1.215035), (23107,-0.979012), (23108,-0.817315), (23109,-0.989585), (23110,-1.061987), (23111,-1.131139), (23112,-0.935999), (23113,-1.085044), (23114,-1.137941), (23115,-0.943720), (23116,-0.919048), (23117,-1.092244), (23118,-1.140031), (23119,-1.330886), (23120,-1.057236), (23121,-1.187703), (23122,-1.233167), (23123,-1.019912), (23124,-0.866568), (23125,-1.023046), (23126,-1.075016), (23127,-1.152064), (23128,-0.959704), (23129,-1.113858), (23130,-1.178834), (23131,-0.942811), (23132,-0.908383), (23133,-1.083445), (23134,-1.107538), (23135,-1.296069), (23136,-0.996872), (23137,-1.126412), (23138,-1.185809), (23139,-0.970230), (23140,-0.826642), (23141,-0.985906), (23142,-1.065277), (23143,-1.111675), (23144,-1.050766), (23145,-1.210963), (23146,-0.848135), (23147,-0.996253), (23148,-0.990622), (23149,-1.139204), (23150,-1.203710), (23151,-1.372729), (23152,-1.112555), (23153,-1.259740), (23154,-0.914101), (23155,-1.051073), (23156,-0.901912), (23157,-1.082541), (23158,-1.055545), (23159,-1.213419), (23160,-0.965787), (23161,-1.097180), (23162,-1.159827), (23163,-0.909408), (23164,-0.891705), (23165,-1.070474), (23166,-1.097823), (23167,-1.299360), (23168,-1.608190), (23169,-1.341980), (23170,-1.083196), (23171,-1.140275), (23172,-1.307435), (23173,-1.143415), (23174,-1.243225), (23175,-1.312377), (23176,-1.480464), (23177,-1.189169), (23178,-0.968481), (23179,-1.001867), (23180,-1.158344), (23181,-1.131348), (23182,-1.286430), (23183,-1.311919), (23184,-1.473506), (23185,-1.231917), (23186,-0.976852), (23187,-0.999086), (23188,-1.187153), (23189,-1.021267), (23190,-1.059769), (23191,-1.120092), (23192,-1.484200), (23193,-1.217527), (23194,-0.955029), (23195,-1.021395), (23196,-1.171836), (23197,-1.149944), (23198,-1.346834), (23199,-1.383939), (23200,-1.561782), (23201,-1.276060), (23202,-1.039574), (23203,-1.079002), (23204,-1.242449), (23205,-1.066813), (23206,-1.153617), (23207,-1.203721), (23208,-1.382497), (23209,-1.106531), (23210,-0.872367), (23211,-0.935947), (23212,-1.088248), (23213,-1.066355), (23214,-1.296689), (23215,-1.356549), (23216,-1.519533), (23217,-1.227311), (23218,-0.990825), (23219,-1.034430), (23220,-1.187657), (23221,-1.040356), (23222,-1.136916), (23223,-1.175411), (23224,-1.581322), (23225,-1.326721), (23226,-1.087448), (23227,-1.128266), (23228,-1.267099), (23229,-1.259608), (23230,-1.456962), (23231,-1.507066), (23232,-1.676085), (23233,-1.375505), (23234,-1.119044), (23235,-1.195629), (23236,-1.355362), (23237,-1.209914), (23238,-1.257239), (23239,-1.318958), (23240,-1.415981), (23241,-1.127936), (23242,-0.902139), (23243,-0.944347), (23244,-1.080856), (23245,-1.066396), (23246,-1.262360), (23247,-1.262302), (23248,-1.445717), (23249,-1.142813), (23250,-0.943020), (23251,-0.987095), (23252,-1.135676), (23253,-0.953072), (23254,-1.034303), (23255,-1.087193), (23256,-1.496361), (23257,-1.262198), (23258,-1.009919), (23259,-1.041915), (23260,-1.203039), (23261,-1.173250), (23262,-1.393828), (23263,-1.427684), (23264,-1.582765), (23265,-1.293330), (23266,-1.034546), (23267,-1.084656), (23268,-1.262499), (23269,-1.125886), (23270,-1.179246), (23271,-1.233070), (23272,-1.277138), (23273,-1.447548), (23274,-0.746571), (23275,-0.890506), (23276,-0.962451), (23277,-1.124038), (23278,-1.152777), (23279,-1.292067), (23280,-1.329635), (23281,-1.484253), (23282,-0.816719), (23283,-0.966697), (23284,-1.048392), (23285,-1.218801), (23286,-0.953981), (23287,-1.070052), (23288,-1.164752), (23289,-0.899005), (23290,-1.070348), (23291,-0.723312), (23292,-0.882576), (23293,-0.871372), (23294,-1.011124), (23295,-1.128122), (23296,-1.239077), (23297,-0.995165), (23298,-1.137704), (23299,-0.798107), (23300,-0.941109), (23301,-0.831434), (23302,-0.941926), (23303,-0.925149), (23304,-1.148051), (23305,-1.287340), (23306,-1.001155), (23307,-0.780930), (23308,-0.827321), (23309,-1.010273), (23310,-0.935432), (23311,-1.141151), (23312,-1.204730), (23313,-1.369567), (23314,-1.077340), (23315,-0.842250), (23316,-0.865886), (23317,-1.034436), (23318,-0.911756), (23319,-0.947001), (23320,-0.859154), (23321,-1.016558), (23322,-1.081071), (23323,-0.847834), (23324,-0.851032), (23325,-0.994968), (23326,-1.046005), (23327,-1.223847), (23328,-0.964606), (23329,-1.129443), (23330,-1.191163), (23331,-0.929599), (23332,-0.753963), (23333,-0.943421), (23334,-0.987489), (23335,-1.043172), (23336,-1.365472), (23337,-1.087182), (23338,-0.853952), (23339,-0.889197), (23340,-1.057747), (23341,-1.035398), (23342,-1.241574), (23343,-1.249882), (23344,-1.416115), (23345,-1.141539), (23346,-0.914345), (23347,-0.983497), (23348,-1.128366), (23349,-0.972236), (23350,-1.073905), (23351,-1.111937), (23352,-0.878237), (23353,-1.035184), (23354,-1.081575), (23355,-0.853911), (23356,-0.840854), (23357,-0.998258), (23358,-1.027931), (23359,-1.230394), (23360,-0.948849), (23361,-1.090931), (23362,-1.141968), (23363,-0.896659), (23364,-0.745175), (23365,-0.910012), (23366,-0.974061), (23367,-1.048786), (23368,-1.194581), (23369,-0.901890), (23370,-1.051405), (23371,-0.712728), (23372,-0.884534), (23373,-0.879366), (23374,-1.034454), (23375,-1.102680), (23376,-1.234999), (23377,-0.989691), (23378,-1.133626), (23379,-0.799602), (23380,-0.924959), (23381,-0.791126), (23382,-0.967579), (23383,-0.928967), (23384,-0.821609), (23385,-1.004568), (23386,-1.043526), (23387,-0.789388), (23388,-0.775398), (23389,-0.957886), (23390,-1.001028), (23391,-1.182589), (23392,-0.906623), (23393,-1.066820), (23394,-1.135973), (23395,-0.869292), (23396,-0.708522), (23397,-0.887298), (23398,-0.941121), (23399,-1.013987), (23400,-1.303312), (23401,-1.004121), (23402,-0.772281), (23403,-0.769900), (23404,-0.969577), (23405,-0.952337), (23406,-1.144581), (23407,-1.164498), (23408,-1.307970), (23409,-1.019925), (23410,-0.753245), (23411,-0.819611), (23412,-0.993277), (23413,-0.855268), (23414,-0.901195), (23415,-0.968488), (23416,-1.395301), (23417,-1.114225), (23418,-0.866593), (23419,-0.919027), (23420,-1.105698), (23421,-1.093561), (23422,-1.261654), (23423,-1.352635), (23424,-1.518868), (23425,-1.259620), (23426,-1.443042), (23427,-1.069068), (23428,-1.227405), (23429,-1.086140), (23430,-1.188736), (23431,-1.158954), (23432,-1.283378), (23433,-1.443575), (23434,-1.150884), (23435,-0.945988), (23436,-1.010031), (23437,-1.154429), (23438,-1.119074), (23439,-1.312245), (23440,-1.369319), (23441,-1.516047), (23442,-1.283743), (23443,-1.010564), (23444,-1.046736), (23445,-1.215755), (23446,-1.073564), (23447,-1.107876), (23448,-1.376763), (23449,-1.526271), (23450,-1.241946), (23451,-1.029617), (23452,-1.051387), (23453,-1.247351), (23454,-1.205027), (23455,-1.395875), (23456,-1.440406), (23457,-1.575519), (23458,-1.317204), (23459,-1.080718), (23460,-1.133152), (23461,-1.276624), (23462,-1.122816), (23463,-1.224022), (23464,-1.452497), (23465,-1.612687), (23466,-0.941441), (23467,-1.118820), (23468,-1.135017), (23469,-1.294281), (23470,-1.298406), (23471,-1.459066), (23472,-1.516609), (23473,-1.660081), (23474,-0.997187), (23475,-1.123471), (23476,-1.213995), (23477,-1.403452), (23478,-1.167429), (23479,-1.319261), (23480,-1.414430), (23481,-1.551860), (23482,-1.275430), (23483,-1.050560), (23484,-1.097877), (23485,-1.256678), (23486,-1.239901), (23487,-1.407525), (23488,-1.454849), (23489,-1.630368), (23490,-1.353012), (23491,-1.105380), (23492,-1.171282), (23493,-1.328686), (23494,-1.177202), (23495,-1.248214), (23496,-1.364285), (23497,-1.501715), (23498,-1.181623), (23499,-0.958605), (23500,-1.002216), (23501,-1.157761), (23502,-1.163745), (23503,-1.326259), (23504,-1.356395), (23505,-1.502190), (23506,-1.237839), (23507,-0.992994), (23508,-1.017550), (23509,-1.185643), (23510,-1.018831), (23511,-1.092629), (23512,-1.417721), (23513,-1.546328), (23514,-1.283367), (23515,-1.018547), (23516,-1.085846), (23517,-1.244646), (23518,-1.219504), (23519,-1.399669), (23520,-1.462785), (23521,-1.599288), (23522,-1.350729), (23523,-1.097061), (23524,-1.130447), (23525,-1.311539), (23526,-1.165171), (23527,-1.262194), (23528,-1.284897), (23529,-1.443697), (23530,-1.171444), (23531,-0.915916), (23532,-0.969277), (23533,-1.115072), (23534,-1.121513), (23535,-1.299362), (23536,-1.322992), (23537,-1.466001), (23538,-1.198394), (23539,-0.958658), (23540,-1.005049), (23541,-1.164319), (23542,-1.023981), (23543,-1.049940), (23544,-1.179474), (23545,-1.358712), (23546,-1.085069), (23547,-0.826285), (23548,-0.881505), (23549,-1.061207), (23550,-1.042571), (23551,-1.245967), (23552,-1.222215), (23553,-1.416782), (23554,-1.132920), (23555,-0.882038), (23556,-0.935399), (23557,-1.084907), (23558,-0.922741), (23559,-1.003045), (23560,-1.212941), (23561,-1.407038), (23562,-1.095306), (23563,-0.843497), (23564,-0.925655), (23565,-1.063554), (23566,-1.049557), (23567,-1.225546), (23568,-1.263115), (23569,-1.427488), (23570,-1.174283), (23571,-0.913176), (23572,-0.973506), (23573,-1.130447), (23574,-0.988255), (23575,-1.056480), (23576,-1.207385), (23577,-0.948607), (23578,-1.074428), (23579,-1.113386), (23580,-0.898271), (23581,-0.852691), (23582,-1.028216), (23583,-1.081107), (23584,-1.251060), (23585,-0.956978), (23586,-1.102767), (23587,-1.177035), (23588,-0.906172), (23589,-0.780706), (23590,-0.914422), (23591,-0.978001), (23592,-1.277546), (23593,-1.045242), (23594,-1.191964), (23595,-0.850037), (23596,-1.011625), (23597,-0.996708), (23598,-1.126241), (23599,-1.176352), (23600,-1.355590), (23601,-1.095416), (23602,-1.216590), (23603,-0.882566), (23604,-1.045080), (23605,-0.889883), (23606,-1.047287), (23607,-1.068600), (23608,-1.365352), (23609,-1.092635), (23610,-1.241687), (23611,-0.928094), (23612,-1.062274), (23613,-1.040851), (23614,-1.214517), (23615,-1.306893), (23616,-1.456402), (23617,-1.172540), (23618,-1.329017), (23619,-1.009388), (23620,-1.144501), (23621,-1.024607), (23622,-1.117447), (23623,-1.065831), (23624,-1.304524), (23625,-1.029021), (23626,-1.201291), (23627,-0.859371), (23628,-0.986581), (23629,-0.978164), (23630,-1.134641), (23631,-1.218659), (23632,-1.397434), (23633,-1.118682), (23634,-1.238929), (23635,-0.943915), (23636,-1.084601), (23637,-0.927544), (23638,-1.114215), (23639,-1.092329), (23640,-1.198174), (23641,-0.884588), (23642,-1.048498), (23643,-1.105108), (23644,-0.880238), (23645,-0.865778), (23646,-1.004140), (23647,-1.089084), (23648,-1.224197), (23649,-0.962163), (23650,-1.144188), (23651,-1.178507), (23652,-0.959209), (23653,-0.791470), (23654,-0.973495), (23655,-1.010600), (23656,-1.448558), (23657,-1.170269), (23658,-0.911955), (23659,-0.969028), (23660,-1.127829), (23661,-1.113375), (23662,-1.300973), (23663,-1.371985), (23664,-1.509415), (23665,-1.219516), (23666,-0.971421), (23667,-1.056365), (23668,-1.193331), (23669,-1.050676), (23670,-1.109609), (23671,-1.164366), (23672,-1.349178), (23673,-1.053237), (23674,-1.202745), (23675,-0.856179), (23676,-0.984786), (23677,-0.993093), (23678,-1.143992), (23679,-1.246124), (23680,-1.608373), (23681,-1.323121), (23682,-1.474952), (23683,-1.131172), (23684,-1.261169), (23685,-1.086467), (23686,-1.248054), (23687,-1.249855), (23688,-1.480653), (23689,-1.210259), (23690,-1.384389), (23691,-1.037353), (23692,-1.176642), (23693,-1.154756), (23694,-1.317269), (23695,-1.385958), (23696,-1.552191), (23697,-1.263683), (23698,-1.407155), (23699,-1.092636), (23700,-1.249114), (23701,-1.140365), (23702,-1.252717), (23703,-1.202960), (23704,-1.467664), (23705,-1.611136), (23706,-1.350499), (23707,-1.103330), (23708,-1.148795), (23709,-1.364263), (23710,-1.312647), (23711,-1.475630), (23712,-1.487645), (23713,-1.662243), (23714,-1.359333), (23715,-1.132139), (23716,-1.179457), (23717,-1.325252), (23718,-1.199786), (23719,-1.286589), (23720,-1.385936), (23721,-1.561918), (23722,-1.262264), (23723,-1.026711), (23724,-1.050341), (23725,-1.240262), (23726,-1.223485), (23727,-1.405510), (23728,-1.463517), (23729,-1.626031), (23730,-1.318481), (23731,-1.111719), (23732,-1.192023), (23733,-1.320166), (23734,-1.127343), (23735,-1.236444), (23736,-1.447730), (23737,-1.633938), (23738,-1.334748), (23739,-1.106157), (23740,-1.189712), (23741,-1.360585), (23742,-1.325230), (23743,-1.504005), (23744,-1.544823), (23745,-1.719416), (23746,-1.454132), (23747,-1.204640), (23748,-1.272402), (23749,-1.414941), (23750,-1.248598), (23751,-1.335402), (23752,-1.407804), (23753,-1.534088), (23754,-1.251159), (23755,-1.011886), (23756,-1.074069), (23757,-1.193390), (23758,-1.204015), (23759,-1.406015), (23760,-1.438937), (23761,-1.599597), (23762,-1.323631), (23763,-1.085748), (23764,-1.139109), (23765,-1.341109), (23766,-1.171046), (23767,-1.217437), (23768,-1.511872), (23769,-1.654881), (23770,-1.361263), (23771,-1.146611), (23772,-1.220409), (23773,-1.370844), (23774,-1.323411), (23775,-1.494753), (23776,-1.552760), (23777,-1.734785), (23778,-1.443954), (23779,-1.202358), (23780,-1.253859), (23781,-1.387581), (23782,-1.244920), (23783,-1.333120), (23784,-1.371152), (23785,-1.517410), (23786,-1.222866), (23787,-0.989166), (23788,-1.059245), (23789,-1.202254), (23790,-1.189660), (23791,-1.357283), (23792,-1.405534), (23793,-1.578730), (23794,-1.276290), (23795,-1.031444), (23796,-1.078768), (23797,-1.225027), (23798,-1.068896), (23799,-1.158487), (23800,-1.264802), (23801,-1.411524), (23802,-1.119766), (23803,-0.866098), (23804,-0.924567), (23805,-1.075935), (23806,-1.050793), (23807,-1.261152), (23808,-1.339597), (23809,-1.491428), (23810,-1.207103), (23811,-0.973866), (23812,-1.038379), (23813,-1.202283), (23814,-1.055451), (23815,-1.113921), (23816,-1.332176), (23817,-1.498403), (23818,-1.217797), (23819,-0.995243), (23820,-1.041640), (23821,-1.212977), (23822,-1.184591), (23823,-1.382872), (23824,-1.417653), (23825,-1.598746), (23826,-1.273081), (23827,-0.997578), (23828,-1.068590), (23829,-1.256188), (23830,-1.121892), (23831,-1.179429), (23832,-1.317791), (23833,-1.072019), (23834,-1.220601), (23835,-1.293003), (23836,-1.034225), (23837,-1.002583), (23838,-1.174389), (23839,-1.235646), (23840,-1.368435), (23841,-1.120803), (23842,-1.259166), (23843,-1.286052), (23844,-1.048169), (23845,-0.889259), (23846,-1.047126), (23847,-1.104669), (23848,-1.444157), (23849,-1.198848), (23850,-1.358575), (23851,-0.972523), (23852,-1.134579), (23853,-1.139167), (23854,-1.278920), (23855,-1.318348), (23856,-1.475752), (23857,-1.210469), (23858,-1.364623), (23859,-1.025489), (23860,-1.162455), (23861,-1.024447), (23862,-1.165132), (23863,-1.151605), (23864,-1.425132), (23865,-1.103644), (23866,-1.266164), (23867,-0.920988), (23868,-1.075605), (23869,-1.058829), (23870,-1.219952), (23871,-1.290031), (23872,-1.442796), (23873,-1.190054), (23874,-1.333990), (23875,-1.011111), (23876,-1.157833), (23877,-0.992417), (23878,-1.146571), (23879,-1.135831), (23880,-1.398212), (23881,-1.128752), (23882,-1.263858), (23883,-0.946552), (23884,-1.107676), (23885,-1.062102), (23886,-1.223219), (23887,-1.288658), (23888,-1.462788), (23889,-1.167780), (23890,-1.325647), (23891,-0.963283), (23892,-1.103042), (23893,-0.984075), (23894,-1.132656), (23895,-1.050382), (23896,-1.186885), (23897,-0.922071), (23898,-1.070653), (23899,-1.156993), (23900,-0.903782), (23901,-0.879109), (23902,-1.036050), (23903,-1.077801), (23904,-1.250534), (23905,-0.991756), (23906,-1.140338), (23907,-1.208557), (23908,-0.967431), (23909,-0.822916), (23910,-0.976144), (23911,-1.002560), (23912,-1.301641), (23913,-1.056326), (23914,-1.221169), (23915,-0.857414), (23916,-1.025038), (23917,-1.025443), (23918,-1.167525), (23919,-1.247823), (23920,-1.388972), (23921,-1.101860), (23922,-1.256941), (23923,-0.928953), (23924,-1.095186), (23925,-0.941849), (23926,-1.094144), (23927,-1.066678), (23928,-1.396416), (23929,-1.124163), (23930,-1.251844), (23931,-0.958689), (23932,-1.103558), (23933,-1.054264), (23934,-1.220034), (23935,-1.278967), (23936,-1.636570), (23937,-1.365250), (23938,-1.503149), (23939,-1.177478), (23940,-1.323273), (23941,-1.197806), (23942,-1.341741), (23943,-1.295234), (23944,-1.445675), (23945,-1.599367), (23946,-1.352198), (23947,-1.074835), (23948,-1.118440), (23949,-1.273064), (23950,-1.279506), (23951,-1.455958), (23952,-1.525574), (23953,-1.683448), (23954,-1.409341), (23955,-1.191897), (23956,-1.240147), (23957,-1.389662), (23958,-1.224239), (23959,-1.298508), (23960,-1.319351), (23961,-1.501376), (23962,-1.207295), (23963,-1.395356), (23964,-1.056216), (23965,-1.204798), (23966,-1.175942), (23967,-1.350072), (23968,-1.452667), (23969,-1.599396), (23970,-1.314137), (23971,-1.455286), (23972,-1.124975), (23973,-1.274020), (23974,-1.093275), (23975,-1.247893), (23976,-1.397871), (23977,-1.564567), (23978,-1.285351), (23979,-1.060944), (23980,-1.076215), (23981,-1.208534), (23982,-1.241457), (23983,-1.427665), (23984,-1.472666), (23985,-1.622174), (23986,-1.352244), (23987,-1.112508), (23988,-1.170515), (23989,-1.303304), (23990,-1.149967), (23991,-1.243734), (23992,-1.544668), (23993,-1.684427), (23994,-1.403814), (23995,-1.171048), (23996,-1.205830), (23997,-1.367880), (23998,-1.372468), (23999,-1.538701), (24000,-1.621786), (24001,-1.781513), (24002,-1.506017), (24003,-1.242586), (24004,-1.267613), (24005,-1.444065), (24006,-1.276789), (24007,-1.345941), (24008,-1.428105), (24009,-1.619417), (24010,-1.310934), (24011,-1.084209), (24012,-1.124558), (24013,-1.256421), (24014,-1.267978), (24015,-1.457899), (24016,-1.487102), (24017,-1.670987), (24018,-1.394094), (24019,-1.162717), (24020,-1.217004), (24021,-1.352117), (24022,-1.182518), (24023,-1.249347), (24024,-1.315713), (24025,-1.455009), (24026,-1.184152), (24027,-1.349452), (24028,-1.001489), (24029,-1.142175), (24030,-1.143050), (24031,-1.324605), (24032,-1.405373), (24033,-1.560454), (24034,-1.269629), (24035,-1.417741), (24036,-1.085107), (24037,-1.218830), (24038,-1.081741), (24039,-1.254017), (24040,-1.217266), (24041,-1.385815), (24042,-1.120532), (24043,-1.240316), (24044,-0.893750), (24045,-1.062300), (24046,-1.066888), (24047,-1.223835), (24048,-1.295310), (24049,-1.437386), (24050,-1.156774), (24051,-1.320684), (24052,-0.972258), (24053,-1.147314), (24054,-0.989330), (24055,-1.152313), (24056,-1.176407), (24057,-1.329634), (24058,-1.060168), (24059,-1.206896), (24060,-0.851500), (24061,-1.006118), (24062,-0.971690), (24063,-1.145819), (24064,-1.223794), (24065,-1.342188), (24066,-1.056466), (24067,-1.228273), (24068,-0.916076), (24069,-1.065121), (24070,-0.893199), (24071,-1.053859), (24072,-1.218696), (24073,-1.327798), (24074,-1.069014), (24075,-1.205053), (24076,-0.888681), (24077,-1.043299), (24078,-1.041851), (24079,-1.180676), (24080,-1.264694), (24081,-1.395624), (24082,-1.115011), (24083,-1.288677), (24084,-0.941641), (24085,-1.079540), (24086,-0.907155), (24087,-1.048304), (24088,-1.395224), (24089,-1.129013), (24090,-1.259017), (24091,-1.280323), (24092,-1.042910), (24093,-1.061901), (24094,-1.199800), (24095,-1.261983), (24096,-1.430069), (24097,-1.184297), (24098,-1.309191), (24099,-1.350009), (24100,-1.105627), (24101,-0.968081), (24102,-1.118522), (24103,-1.188138), (24104,-1.273082), (24105,-0.994330), (24106,-1.158703), (24107,-1.201844), (24108,-0.943530), (24109,-0.935113), (24110,-1.120388), (24111,-1.180717), (24112,-1.359956), (24113,-1.057509), (24114,-1.204237), (24115,-1.261774), (24116,-1.042476), (24117,-0.891925), (24118,-1.048866), (24119,-1.118482), (24120,-1.320018), (24121,-1.017108), (24122,-1.192170), (24123,-1.244134), (24124,-0.995575), (24125,-0.978329), (24126,-1.132484), (24127,-1.210928), (24128,-1.366942), (24129,-1.057996), (24130,-1.218656), (24131,-1.275266), (24132,-1.015556), (24133,-0.887302), (24134,-1.043780), (24135,-1.093421), (24136,-1.274056), (24137,-0.999943), (24138,-1.161530), (24139,-1.184233), (24140,-0.979337), (24141,-0.964414), (24142,-1.099990), (24143,-1.161247), (24144,-1.341882), (24145,-1.065446), (24146,-1.223320), (24147,-1.260888), (24148,-1.049023), (24149,-0.891966), (24150,-1.034042), (24151,-1.097158), (24152,-1.364648), (24153,-1.066854), (24154,-1.251666), (24155,-1.336146), (24156,-1.072722), (24157,-1.052226), (24158,-1.231465), (24159,-1.274606), (24160,-1.444089), (24161,-1.149075), (24162,-1.288834), (24163,-1.372852), (24164,-1.100135), (24165,-0.952834), (24166,-1.131140), (24167,-1.166855), (24168,-1.355379), (24169,-1.113784), (24170,-1.243324), (24171,-0.892574), (24172,-1.054161), (24173,-1.040171), (24174,-1.183173), (24175,-1.251862), (24176,-1.432961), (24177,-1.152812), (24178,-1.289784), (24179,-0.961790), (24180,-1.095043), (24181,-0.967253), (24182,-1.095860), (24183,-1.091162), (24184,-1.458984), (24185,-1.156537), (24186,-1.325556), (24187,-1.024512), (24188,-1.142437), (24189,-1.131233), (24190,-1.268199), (24191,-1.351753), (24192,-1.423229), (24193,-1.570414), (24194,-1.325105), (24195,-1.050529), (24196,-1.119218), (24197,-1.267336), (24198,-1.100530), (24199,-1.205449), (24200,-1.376785), (24201,-1.534196), (24202,-1.240578), (24203,-0.990623), (24204,-1.054202), (24205,-1.206033), (24206,-1.217591), (24207,-1.397756), (24208,-1.459476), (24209,-1.596448), (24210,-1.299111), (24211,-1.110470), (24212,-1.142929), (24213,-1.323095), (24214,-1.145606), (24215,-1.221721), (24216,-1.459488), (24217,-1.517494), (24218,-1.669789), (24219,-1.007828), (24220,-1.183354), (24221,-1.255293), (24222,-1.387149), (24223,-1.370836), (24224,-1.529173), (24225,-1.560236), (24226,-1.698598), (24227,-1.043143), (24228,-1.204261), (24229,-1.231610), (24230,-1.407136), (24231,-1.167863), (24232,-1.345705), (24233,-1.417181), (24234,-1.577841), (24235,-0.897765), (24236,-1.046810), (24237,-1.086232), (24238,-1.267331), (24239,-1.270992), (24240,-1.452084), (24241,-1.473861), (24242,-1.637771), (24243,-0.938647), (24244,-1.098844), (24245,-1.150345), (24246,-1.308218), (24247,-1.075445), (24248,-1.360594), (24249,-1.413948), (24250,-1.563926), (24251,-0.875491), (24252,-1.058906), (24253,-1.135491), (24254,-1.329595), (24255,-1.349048), (24256,-1.483691), (24257,-1.544484), (24258,-1.682384), (24259,-0.982797), (24260,-1.162035), (24261,-1.198671), (24262,-1.376056), (24263,-1.137710), (24264,-1.324845), (24265,-1.387497), (24266,-1.560693), (24267,-0.866686), (24268,-1.006902), (24269,-1.066768), (24270,-1.215813), (24271,-1.262667), (24272,-1.401499), (24273,-1.450213), (24274,-1.620160), (24275,-0.934511), (24276,-1.073800), (24277,-1.158281), (24278,-1.285035), (24279,-1.079206), (24280,-1.462819), (24281,-1.540800), (24282,-1.670797), (24283,-0.983759), (24284,-1.141626), (24285,-1.208925), (24286,-1.351001), (24287,-1.403434), (24288,-1.551083), (24289,-1.635564), (24290,-1.733983), (24291,-1.064126), (24292,-1.221067), (24293,-1.238661), (24294,-1.383060), (24295,-1.169804), (24296,-1.335104), (24297,-1.374063), (24298,-1.525901), (24299,-0.861147), (24300,-1.040849), (24301,-1.074241), (24302,-1.197275), (24303,-1.219515), (24304,-1.362987), (24305,-1.417274), (24306,-1.597439), (24307,-0.886707), (24308,-1.085457), (24309,-1.139744), (24310,-1.284142), (24311,-1.043943), (24312,-1.222718), (24313,-1.283511), (24314,-1.429306), (24315,-0.773382), (24316,-0.910812), (24317,-0.983683), (24318,-1.167098), (24319,-1.171687), (24320,-1.291007), (24321,-1.371312), (24322,-1.514314), (24323,-0.833775), (24324,-0.979107), (24325,-1.036644), (24326,-1.201487), (24327,-0.989615), (24328,-1.298915), (24329,-1.395005), (24330,-1.534301), (24331,-0.833324), (24332,-1.010703), (24333,-1.047801), (24334,-1.176414), (24335,-1.208867), (24336,-1.375563), (24337,-1.439613), (24338,-1.576115), (24339,-0.890467), (24340,-1.074345), (24341,-1.137925), (24342,-1.312517), (24343,-1.024942), (24344,-1.141470), (24345,-1.281692), (24346,-1.019195), (24347,-1.214226), (24348,-0.860690), (24349,-1.021350), (24350,-0.980880), (24351,-1.113669), (24352,-1.193504), (24353,-1.341159), (24354,-1.063333), (24355,-1.225847), (24356,-0.920156), (24357,-1.060842), (24358,-0.944198), (24359,-1.071872), (24360,-1.295706), (24361,-1.461933), (24362,-1.194333), (24363,-0.944841), (24364,-0.979153), (24365,-1.154215), (24366,-1.127213), (24367,-1.326890), (24368,-1.386756), (24369,-1.553453), (24370,-1.243110), (24371,-0.995942), (24372,-0.999603), (24373,-1.186738), (24374,-1.035723), (24375,-1.135063), (24376,-1.286431), (24377,-1.441982), (24378,-1.160906), (24379,-0.922097), (24380,-1.027485), (24381,-1.159342), (24382,-1.145352), (24383,-1.315298), (24384,-1.372841), (24385,-1.533965), (24386,-1.251956), (24387,-1.007574), (24388,-1.068830), (24389,-1.198834), (24390,-1.048746), (24391,-1.116508), (24392,-1.273912), (24393,-1.459657), (24394,-1.209702), (24395,-0.937912), (24396,-0.991736), (24397,-1.122666), (24398,-1.144442), (24399,-1.335760), (24400,-1.379365), (24401,-1.504258), (24402,-1.223646), (24403,-0.965795), (24404,-1.044703), (24405,-1.204893), (24406,-1.023222), (24407,-1.126744), (24408,-1.153167), (24409,-1.314754), (24410,-1.018813), (24411,-1.149743), (24412,-0.798061), (24413,-0.960118), (24414,-0.950304), (24415,-1.105391), (24416,-1.207518), (24417,-1.375611), (24418,-1.094535), (24419,-1.245440), (24420,-0.921165), (24421,-1.065100), (24422,-0.941956), (24423,-1.071490), (24424,-1.265131), (24425,-1.435077), (24426,-1.149355), (24427,-0.892900), (24428,-0.957870), (24429,-1.105988), (24430,-1.099430), (24431,-1.294924), (24432,-1.350138), (24433,-1.491757), (24434,-1.184201), (24435,-0.968622), (24436,-1.000148), (24437,-1.174740), (24438,-0.994459), (24439,-1.078946), (24440,-1.269794), (24441,-1.397937), (24442,-1.109429), (24443,-0.894314), (24444,-0.935132), (24445,-1.093463), (24446,-1.095265), (24447,-1.290765), (24448,-1.277702), (24449,-1.427210), (24450,-0.749457), (24451,-0.895716), (24452,-0.973227), (24453,-1.103694), (24454,-0.851879), (24455,-1.008826), (24456,-1.064040), (24457,-1.219591), (24458,-0.520474), (24459,-0.688560), (24460,-0.765145), (24461,-0.916976), (24462,-0.920174), (24463,-1.071542), (24464,-1.144408), (24465,-1.293459), (24466,-0.626852), (24467,-0.801445), (24468,-0.861768), (24469,-0.986662), (24470,-0.774796), (24471,-0.912696), (24472,-1.181113), (24473,-1.242839), (24474,-1.017498), (24475,-0.716448), (24476,-0.882681), (24477,-0.952303), (24478,-1.178918), (24479,-1.139380), (24480,-1.281456), (24481,-1.325993), (24482,-1.052814), (24483,-0.790780), (24484,-0.954226), (24485,-1.011300), (24486,-1.082312), (24487,-0.944766), (24488,-1.148156), (24489,-1.190371), (24490,-0.949702), (24491,-0.634256), (24492,-0.802343), (24493,-0.843167), (24494,-1.019613), (24495,-0.985185), (24496,-1.149558), (24497,-1.199205), (24498,-0.959469), (24499,-0.679784), (24500,-0.845554), (24501,-0.893804), (24502,-0.930440), (24503,-0.793827), (24504,-1.182550), (24505,-1.247056), (24506,-1.027295), (24507,-0.709526), (24508,-0.852065), (24509,-0.917504), (24510,-1.129723), (24511,-1.121769), (24512,-1.276850), (24513,-1.314882), (24514,-1.085365), (24515,-0.814972), (24516,-0.983065), (24517,-1.053144), (24518,-1.119509), (24519,-0.971745), (24520,-1.052512), (24521,-1.105409), (24522,-0.905153), (24523,-0.590634), (24524,-0.754081), (24525,-0.819050), (24526,-0.969955), (24527,-0.975939), (24528,-1.125911), (24529,-1.171375), (24530,-0.937676), (24531,-0.635698), (24532,-0.811224), (24533,-0.850646), (24534,-0.899360), (24535,-0.754382), (24536,-1.164013), (24537,-1.212263), (24538,-0.980887), (24539,-0.709097), (24540,-0.854429), (24541,-0.894784), (24542,-1.074949), (24543,-1.074897), (24544,-1.226265), (24545,-1.262901), (24546,-1.005976), (24547,-0.736516), (24548,-0.892067), (24549,-0.942171), (24550,-1.017366), (24551,-0.861699), (24552,-1.059053), (24553,-1.122169), (24554,-0.910304), (24555,-0.593461), (24556,-0.740646), (24557,-0.799586), (24558,-0.989507), (24559,-0.957395), (24560,-1.159859), (24561,-1.181635), (24562,-0.989745), (24563,-0.684511), (24564,-0.813582), (24565,-0.868338), (24566,-0.932844), (24567,-0.795299), (24568,-0.836580), (24569,-0.896447), (24570,-1.017621), (24571,-0.348228), (24572,-0.503778), (24573,-0.578967), (24574,-0.723372), (24575,-0.743289), (24576,-0.925777), (24577,-0.980991), (24578,-1.120750), (24579,-0.426736), (24580,-0.600865), (24581,-0.654225), (24582,-0.791198), (24583,-0.575613), (24584,-0.892809), (24585,-0.950345), (24586,-1.058521), (24587,-0.351964), (24588,-0.511692), (24589,-0.583637), (24590,-0.757759), (24591,-0.778146), (24592,-0.905356), (24593,-0.976832), (24594,-1.109621), (24595,-0.451843), (24596,-0.586023), (24597,-0.653785), (24598,-0.795398), (24599,-0.581673), (24600,-0.863565), (24601,-1.035835), (24602,-0.751973), (24603,-0.503407), (24604,-0.569773), (24605,-0.714642), (24606,-0.700651), (24607,-0.897536), (24608,-0.936037), (24609,-1.126421), (24610,-0.824908), (24611,-0.579599), (24612,-0.645965), (24613,-0.799656), (24614,-0.681152), (24615,-0.765169), (24616,-1.085145), (24617,-1.218398), (24618,-0.536000), (24619,-0.676222), (24620,-0.726332), (24621,-0.871194), (24622,-0.879965), (24623,-1.037839), (24624,-1.084230), (24625,-1.235598), (24626,-0.562022), (24627,-0.724073), (24628,-0.776970), (24629,-0.898614), (24630,-0.683956), (24631,-0.819532), (24632,-0.830162), (24633,-0.993603), (24634,-0.720423), (24635,-0.469078), (24636,-0.523365), (24637,-0.681239), (24638,-0.686754), (24639,-0.881321), (24640,-0.947687), (24641,-1.112524), (24642,-0.824022), (24643,-0.591249), (24644,-0.629744), (24645,-0.783905), (24646,-0.615695), (24647,-0.685781), (24648,-0.847368), (24649,-1.002919), (24650,-0.723696), (24651,-0.476064), (24652,-0.515029), (24653,-0.650136), (24654,-0.658443), (24655,-0.828390), (24656,-0.878500), (24657,-1.039624), (24658,-0.798955), (24659,-0.542963), (24660,-0.580068), (24661,-0.769990), (24662,-0.624078), (24663,-0.737826), (24664,-0.881298), (24665,-1.017801), (24666,-0.744621), (24667,-0.499776), (24668,-0.547094), (24669,-0.716113), (24670,-0.692367), (24671,-0.853028), (24672,-0.893846), (24673,-1.054970), (24674,-0.787363), (24675,-0.553669), (24676,-0.617249), (24677,-0.775116), (24678,-0.635711), (24679,-0.723442), (24680,-0.981183), (24681,-1.112113), (24682,-0.439933), (24683,-0.580155), (24684,-0.660453), (24685,-0.810431), (24686,-0.818269), (24687,-0.972424), (24688,-1.029034), (24689,-1.183188), (24690,-0.495680), (24691,-0.625220), (24692,-0.701805), (24693,-0.839241), (24694,-0.618083), (24695,-0.750403), (24696,-1.038801), (24697,-1.177627), (24698,-0.525422), (24699,-0.703728), (24700,-0.746869), (24701,-0.901487), (24702,-0.913508), (24703,-1.055590), (24704,-1.099658), (24705,-1.255209), (24706,-0.725626), (24707,-0.869098), (24708,-0.913636), (24709,-1.068717), (24710,-0.686384), (24711,-0.861440), (24712,-1.058793), (24713,-1.184150), (24714,-0.775337), (24715,-0.949002), (24716,-0.986108), (24717,-1.163486), (24718,-0.903776), (24719,-1.045851), (24720,-1.116400), (24721,-1.282633), (24722,-0.729363), (24723,-0.883980), (24724,-0.935487), (24725,-1.079423), (24726,-0.719845), (24727,-0.891651), (24728,-0.903208), (24729,-1.072691), (24730,-1.048945), (24731,-0.805026), (24732,-0.864429), (24733,-1.038095), (24734,-0.770019), (24735,-0.937648), (24736,-0.991008), (24737,-1.131694), (24738,-0.988106), (24739,-0.750230), (24740,-0.811486), (24741,-0.973536), (24742,-0.673882), (24743,-0.730492), (24744,-0.946888), (24745,-0.984920), (24746,-0.780487), (24747,-0.797154), (24748,-0.936443), (24749,-0.977261), (24750,-1.152323), (24751,-0.882857), (24752,-1.046767), (24753,-1.096878), (24754,-0.862714), (24755,-0.698225), (24756,-0.849130), (24757,-0.870906), (24758,-0.939595), (24759,-0.683597), (24760,-1.083936), (24761,-1.246456), (24762,-0.827423), (24763,-0.970895), (24764,-1.000098), (24765,-1.154722), (24766,-0.904767), (24767,-1.061708), (24768,-1.109958), (24769,-1.258540), (24770,-0.728957), (24771,-0.871039), (24772,-0.924863), (24773,-1.111998), (24774,-0.749633), (24775,-0.893105), (24776,-1.008706), (24777,-1.076005), (24778,-0.817221), (24779,-0.792548), (24780,-0.966214), (24781,-1.067883), (24782,-1.212282), (24783,-0.942816), (24784,-1.097440), (24785,-1.157763), (24786,-0.940325), (24787,-0.778622), (24788,-0.933709), (24789,-1.001465), (24790,-1.029747), (24791,-0.752848), (24792,-0.889351), (24793,-1.063480), (24794,-1.045314), (24795,-0.816723), (24796,-0.874730), (24797,-1.042353), (24798,-0.767314), (24799,-0.956308), (24800,-1.015705), (24801,-1.154537), (24802,-0.975645), (24803,-0.740092), (24804,-0.769295), (24805,-0.947607), (24806,-0.656312), (24807,-0.700844), (24808,-0.792294), (24809,-0.835435), (24810,-0.975657), (24811,-0.580782), (24812,-0.746082), (24813,-0.768785), (24814,-0.902038), (24815,-0.665089), (24816,-0.847577), (24817,-0.880036), (24818,-1.036983), (24819,-0.492072), (24820,-0.639727), (24821,-0.726994), (24822,-0.880216), (24823,-0.523893), (24824,-0.704992), (24825,-0.821057), (24826,-0.815889), (24827,-0.566404), (24828,-0.617441), (24829,-0.771595), (24830,-0.529073), (24831,-0.749651), (24832,-0.754703), (24833,-0.925576), (24834,-0.805218), (24835,-0.562233), (24836,-0.605374), (24837,-0.772070), (24838,-0.500281), (24839,-0.579189), (24840,-0.771896), (24841,-0.808075), (24842,-0.981271), (24843,-0.563634), (24844,-0.731727), (24845,-0.779045), (24846,-0.908585), (24847,-0.660020), (24848,-0.820680), (24849,-0.874041), (24850,-1.020299), (24851,-0.476784), (24852,-0.628616), (24853,-0.692195), (24854,-0.868647), (24855,-0.473302), (24856,-0.833697), (24857,-0.971597), (24858,-0.979435), (24859,-0.757350), (24860,-0.842294), (24861,-0.976474), (24862,-0.713050), (24863,-0.890899), (24864,-0.931717), (24865,-1.088194), (24866,-0.906053), (24867,-0.643093), (24868,-0.713641), (24869,-0.880338), (24870,-0.595543), (24871,-0.686993), (24872,-0.727811), (24873,-0.882899), (24874,-0.856360), (24875,-0.606874), (24876,-0.662558), (24877,-0.817176), (24878,-0.525881), (24879,-0.738100), (24880,-0.787277), (24881,-0.962797), (24882,-0.842439), (24883,-0.611526), (24884,-0.645845), (24885,-0.774915), (24886,-0.518460), (24887,-0.602478), (24888,-0.745950), (24889,-0.924719), (24890,-0.946495), (24891,-0.674242), (24892,-0.721103), (24893,-0.882227), (24894,-0.618796), (24895,-0.803145), (24896,-0.842109), (24897,-0.997190), (24898,-0.852676), (24899,-0.627342), (24900,-0.676519), (24901,-0.837179), (24902,-0.554707), (24903,-0.642908), (24904,-0.771514), (24905,-0.903371), (24906,-0.910282), (24907,-0.667296), (24908,-0.722053), (24909,-0.858093), (24910,-0.603955), (24911,-0.803168), (24912,-0.816579), (24913,-0.996751), (24914,-0.839230), (24915,-0.589739), (24916,-0.610119), (24917,-0.761023), (24918,-0.505026), (24919,-0.570928), (24920,-0.821237), (24921,-1.004189), (24922,-1.038044), (24923,-0.793198), (24924,-0.792677), (24925,-0.961697), (24926,-0.667146), (24927,-0.850567), (24928,-0.915537), (24929,-1.038107), (24930,-0.908921), (24931,-0.649680), (24932,-0.701644), (24933,-0.861835), (24934,-0.594234), (24935,-0.668496), (24936,-0.852844), (24937,-1.015358), (24938,-0.591216), (24939,-0.755126), (24940,-0.784798), (24941,-0.939886), (24942,-0.690857), (24943,-0.814355), (24944,-0.903482), (24945,-1.016760), (24946,-0.471385), (24947,-0.613467), (24948,-0.689589), (24949,-0.824695), (24950,-0.476269), (24951,-0.640179), (24952,-0.920675), (24953,-1.066471), (24954,-0.686461), (24955,-0.840152), (24956,-0.893512), (24957,-1.060672), (24958,-0.793065), (24959,-0.964871), (24960,-1.150146), (24961,-1.278290), (24962,-0.704587), (24963,-0.881503), (24964,-0.919998), (24965,-1.096914), (24966,-0.731763), (24967,-0.928190), (24968,-1.047504), (24969,-1.086932), (24970,-0.848586), (24971,-0.835059), (24972,-0.985501), (24973,-1.029569), (24974,-1.246897), (24975,-0.935164), (24976,-1.088855), (24977,-1.140819), (24978,-0.925241), (24979,-0.769111), (24980,-0.923735), (24981,-0.985454), (24982,-1.046711), (24983,-0.738691), (24984,-0.885419), (24985,-0.948066), (24986,-1.092001), (24987,-0.704095), (24988,-0.848030), (24989,-0.869343), (24990,-1.053685), (24991,-0.828815), (24992,-0.990865), (24993,-1.050731), (24994,-1.207672), (24995,-0.646506), (24996,-0.805306), (24997,-0.828942), (24998,-0.986810), (24999,-0.617482), (25000,-1.028040), (25001,-1.093009), (25002,-0.818903), (25003,-0.825344), (25004,-0.979505), (25005,-1.048657), (25006,-1.230683), (25007,-0.961679), (25008,-1.113047), (25009,-1.149226), (25010,-0.933641), (25011,-0.785413), (25012,-0.957219), (25013,-0.985032), (25014,-1.059294), (25015,-0.797260), (25016,-1.148826), (25017,-1.188254), (25018,-0.965700), (25019,-0.905261), (25020,-1.070561), (25021,-1.101630), (25022,-1.269253), (25023,-1.016048), (25024,-1.167879), (25025,-1.224959), (25026,-1.000552), (25027,-0.834666), (25028,-0.988357), (25029,-1.009670), (25030,-1.076962), (25031,-0.747115), (25032,-0.959334), (25033,-1.018730), (25034,-0.805005), (25035,-0.785442), (25036,-0.925195), (25037,-0.969269), (25038,-1.128069), (25039,-0.848384), (25040,-1.002075), (25041,-1.035930), (25042,-0.845430), (25043,-0.693482), (25044,-0.832772), (25045,-0.910753), (25046,-0.985478), (25047,-0.675141), (25048,-0.835332), (25049,-0.943038), (25050,-1.123673), (25051,-0.695817), (25052,-0.833710), (25053,-0.898686), (25054,-1.046334), (25055,-0.801025), (25056,-0.968655), (25057,-1.028978), (25058,-1.172450), (25059,-0.647514), (25060,-0.802138), (25061,-0.859675), (25062,-0.992464), (25063,-0.638929), (25064,-0.785651), (25065,-0.866418), (25066,-1.010354), (25067,-0.596900), (25068,-0.779388), (25069,-0.816957), (25070,-0.972965), (25071,-0.746234), (25072,-0.861842), (25073,-0.906373), (25074,-1.040089), (25075,-0.509580), (25076,-0.663271), (25077,-0.722204), (25078,-0.837342), (25079,-0.481947), (25080,-0.687666), (25081,-0.729411), (25082,-0.885889), (25083,-0.488690), (25084,-0.680008), (25085,-0.744051), (25086,-0.894022), (25087,-0.655219), (25088,-0.832598), (25089,-0.880849), (25090,-1.016425), (25091,-0.477550), (25092,-0.612200), (25093,-0.659524), (25094,-0.821574), (25095,-0.459209), (25096,-0.779655), (25097,-0.827442), (25098,-0.984383), (25099,-0.583002), (25100,-0.716255), (25101,-0.764043), (25102,-0.925630), (25103,-0.673815), (25104,-0.841908), (25105,-0.916633), (25106,-1.053136), (25107,-0.507767), (25108,-0.671208), (25109,-0.752439), (25110,-0.854108), (25111,-0.494993), (25112,-0.862358), (25113,-1.010470), (25114,-0.995553), (25115,-0.782754), (25116,-0.804531), (25117,-0.972154), (25118,-0.693865), (25119,-0.885182), (25120,-0.926464), (25121,-1.065290), (25122,-0.919385), (25123,-0.694977), (25124,-0.740442), (25125,-0.906205), (25126,-0.627453), (25127,-0.684996), (25128,-0.763441), (25129,-0.916662), (25130,-0.903135), (25131,-0.663399), (25132,-0.697254), (25133,-0.833757), (25134,-0.568937), (25135,-0.726347), (25136,-0.818261), (25137,-0.981238), (25138,-0.825114), (25139,-0.553324), (25140,-0.627586), (25141,-0.771528), (25142,-0.502988), (25143,-0.575396), (25144,-0.761598), (25145,-0.887418), (25146,-0.861819), (25147,-0.625333), (25148,-0.686126), (25149,-0.854682), (25150,-0.571283), (25151,-0.735194), (25152,-0.795517), (25153,-0.951531), (25154,-0.802370), (25155,-0.542196), (25156,-0.609495), (25157,-0.773405), (25158,-0.488610), (25159,-0.578200), (25160,-0.689162), (25161,-0.839596), (25162,-0.847441), (25163,-0.624423), (25164,-0.634584), (25165,-0.761338), (25166,-0.517882), (25167,-0.690621), (25168,-0.763023), (25169,-0.894886), (25170,-0.746652), (25171,-0.521318), (25172,-0.583964), (25173,-0.733479), (25174,-0.472841), (25175,-0.511800), (25176,-0.753279), (25177,-0.907897), (25178,-0.899017), (25179,-0.644885), (25180,-0.706605), (25181,-0.855650), (25182,-0.601048), (25183,-0.790043), (25184,-0.846189), (25185,-0.976656), (25186,-0.842360), (25187,-0.599374), (25188,-0.633687), (25189,-0.812925), (25190,-0.510485), (25191,-0.587996), (25192,-0.868493), (25193,-0.917677), (25194,-0.673294), (25195,-0.699247), (25196,-0.834823), (25197,-0.859386), (25198,-1.061849), (25199,-0.786810), (25200,-0.928892), (25201,-0.976673), (25202,-0.730438), (25203,-0.630512), (25204,-0.777234), (25205,-0.790651), (25206,-0.863053), (25207,-0.608922), (25208,-0.933080), (25209,-1.049608), (25210,-0.645441), (25211,-0.775444), (25212,-0.829737), (25213,-1.024298), (25214,-0.746479), (25215,-0.898774), (25216,-0.983254), (25217,-1.014787), (25218,-1.207494), (25219,-0.656547), (25220,-0.816737), (25221,-0.872884), (25222,-1.019143), (25223,-0.685118), (25224,-0.934494), (25225,-0.971129), (25226,-1.114601), (25227,-0.702538), (25228,-0.858552), (25229,-0.916095), (25230,-1.086968), (25231,-0.852811), (25232,-0.991174), (25233,-1.063113), (25234,-1.153630), (25235,-0.618474), (25236,-0.787030), (25237,-0.864079), (25238,-1.000118), (25239,-0.637296), (25240,-0.921042), (25241,-0.996237), (25242,-1.118338), (25243,-0.725323), (25244,-0.865075), (25245,-0.944446), (25246,-1.078632), (25247,-0.849115), (25248,-0.999087), (25249,-1.049198), (25250,-1.201029), (25251,-0.633363), (25252,-0.847899), (25253,-0.874321), (25254,-1.021970), (25255,-0.628491), (25256,-0.961942), (25257,-1.119810), (25258,-0.751872), (25259,-0.911606), (25260,-0.884604), (25261,-1.069415), (25262,-1.119526), (25263,-1.266717), (25264,-0.999574), (25265,-1.143973), (25266,-0.813662), (25267,-0.979895), (25268,-0.837240), (25269,-1.007186), (25270,-0.987623), (25271,-1.123193), (25272,-0.982861), (25273,-1.042257), (25274,-1.193162), (25275,-0.775989), (25276,-0.950118), (25277,-0.996979), (25278,-1.143237), (25279,-0.922080), (25280,-1.055333), (25281,-1.160252), (25282,-1.289791), (25283,-0.760209), (25284,-0.888816), (25285,-0.969120), (25286,-1.132560), (25287,-0.755800), (25288,-0.833312), (25289,-1.000478), (25290,-1.011102), (25291,-0.779726), (25292,-0.780137), (25293,-0.946834), (25294,-0.974647), (25295,-1.142270), (25296,-0.850975), (25297,-1.004666), (25298,-1.026443), (25299,-0.783920), (25300,-0.657057), (25301,-0.779621), (25302,-0.843670), (25303,-0.930005), (25304,-0.963860), (25305,-1.033475), (25306,-1.176021), (25307,-0.715185), (25308,-0.904173), (25309,-0.950101), (25310,-1.129340), (25311,-0.844087), (25312,-1.043764), (25313,-1.093405), (25314,-1.254065), (25315,-0.680357), (25316,-0.830328), (25317,-0.911096), (25318,-1.070360), (25319,-0.714501), (25320,-0.716766), (25321,-0.896468), (25322,-0.917782), (25323,-0.665503), (25324,-0.672878), (25325,-0.824246), (25326,-0.876680), (25327,-1.081460), (25328,-0.815713), (25329,-0.952685), (25330,-1.012545), (25331,-0.776065), (25332,-0.632940), (25333,-0.767126), (25334,-0.813517), (25335,-0.898461), (25336,-0.852887), (25337,-0.882090), (25338,-1.021379), (25339,-0.646942), (25340,-0.810852), (25341,-0.864676), (25342,-1.019300), (25343,-0.755407), (25344,-0.895629), (25345,-0.944806), (25346,-1.071560), (25347,-0.521539), (25348,-0.670121), (25349,-0.757851), (25350,-0.909689), (25351,-0.541751), (25352,-0.730276), (25353,-0.900692), (25354,-0.945693), (25355,-0.736608), (25356,-0.734233), (25357,-0.838689), (25358,-0.917127), (25359,-1.105658), (25360,-0.817150), (25361,-0.966658), (25362,-1.037670), (25363,-0.797471), (25364,-0.632054), (25365,-0.793641), (25366,-0.852575), (25367,-0.898966), (25368,-0.816692), (25369,-0.884917), (25370,-1.052547), (25371,-0.657202), (25372,-0.806247), (25373,-0.840102), (25374,-0.975209), (25375,-0.728510), (25376,-0.919821), (25377,-0.962962), (25378,-1.119903), (25379,-0.637702), (25380,-0.782571), (25381,-0.821066), (25382,-0.959892), (25383,-0.590101), (25384,-0.818575), (25385,-0.886794), (25386,-1.044205), (25387,-0.649323), (25388,-0.766784), (25389,-0.789024), (25390,-0.912058), (25391,-0.661176), (25392,-0.825086), (25393,-0.877514), (25394,-1.040497), (25395,-0.462142), (25396,-0.597255), (25397,-0.676626), (25398,-0.847969), (25399,-0.473069), (25400,-0.829738), (25401,-0.904933), (25402,-1.055374), (25403,-0.660956), (25404,-0.821616), (25405,-0.870330), (25406,-1.004047), (25407,-0.757348), (25408,-0.901283), (25409,-0.972295), (25410,-1.132023), (25411,-0.593617), (25412,-0.738486), (25413,-0.798346), (25414,-0.961792), (25415,-0.602677), (25416,-0.842767), (25417,-0.916102), (25418,-1.064214), (25419,-0.676771), (25420,-0.827213), (25421,-0.881500), (25422,-1.013363), (25423,-0.783376), (25424,-0.921275), (25425,-0.992287), (25426,-1.133899), (25427,-0.548118), (25428,-0.731534), (25429,-0.782571), (25430,-0.934872), (25431,-0.553002), (25432,-0.783799), (25433,-0.847372), (25434,-0.996887), (25435,-0.599219), (25436,-0.781244), (25437,-0.849006), (25438,-0.986442), (25439,-0.743450), (25440,-0.890642), (25441,-0.945392), (25442,-1.111162), (25443,-0.549532), (25444,-0.703686), (25445,-0.790954), (25446,-0.940462), (25447,-0.570671), (25448,-0.926414), (25449,-0.988603), (25450,-0.741898), (25451,-0.745559), (25452,-0.874629), (25453,-0.901052), (25454,-1.103979), (25455,-0.843804), (25456,-0.979380), (25457,-1.001151), (25458,-0.784176), (25459,-0.671714), (25460,-0.823082), (25461,-0.881552), (25462,-0.936303), (25463,-0.652904), (25464,-0.867909), (25465,-0.933812), (25466,-1.068461), (25467,-0.609479), (25468,-0.784541), (25469,-0.855547), (25470,-0.994842), (25471,-0.732345), (25472,-1.069973), (25473,-1.108938), (25474,-1.265878), (25475,-0.729796), (25476,-0.883024), (25477,-0.933128), (25478,-1.060808), (25479,-0.706809), (25480,-0.880475), (25481,-0.981211), (25482,-1.115854), (25483,-0.710297), (25484,-0.879316), (25485,-0.920598), (25486,-1.064533), (25487,-0.802506), (25488,-0.947831), (25489,-1.000728), (25490,-1.162315), (25491,-0.603472), (25492,-0.755773), (25493,-0.801700), (25494,-0.970250), (25495,-0.599533), (25496,-0.964104), (25497,-1.006776), (25498,-1.153504), (25499,-0.772098), (25500,-0.913710), (25501,-0.964284), (25502,-1.139803), (25503,-0.881489), (25504,-1.027284), (25505,-1.074602), (25506,-1.212501), (25507,-0.662486), (25508,-0.793880), (25509,-0.883933), (25510,-1.077104), (25511,-0.685015), (25512,-0.802013), (25513,-0.963600), (25514,-1.018357), (25515,-0.778621), (25516,-0.745583), (25517,-0.913206), (25518,-0.942415), (25519,-1.129086), (25520,-0.833145), (25521,-1.014707), (25522,-1.058775), (25523,-0.804174), (25524,-0.655946), (25525,-0.826356), (25526,-0.854632), (25527,-0.940972), (25528,-0.952066), (25529,-1.082533), (25530,-1.120565), (25531,-0.853421), (25532,-0.833395), (25533,-1.018670), (25534,-1.052982), (25535,-1.231757), (25536,-0.974833), (25537,-1.149895), (25538,-1.157270), (25539,-0.957477), (25540,-0.792524), (25541,-1.006603), (25542,-1.036739), (25543,-1.091026), (25544,-0.765824), (25545,-0.916265), (25546,-1.007246), (25547,-0.780515), (25548,-0.774884), (25549,-0.975024), (25550,-1.007020), (25551,-1.191368), (25552,-0.868953), (25553,-1.020784), (25554,-1.085290), (25555,-0.824653), (25556,-0.682924), (25557,-0.860773), (25558,-0.889513), (25559,-0.956342), (25560,-0.920054), (25561,-1.087220), (25562,-1.141044), (25563,-0.893412), (25564,-0.873379), (25565,-1.017778), (25566,-1.097619), (25567,-1.262455), (25568,-0.965124), (25569,-1.120206), (25570,-1.156847), (25571,-0.909209), (25572,-0.752622), (25573,-0.923031), (25574,-0.961526), (25575,-1.070165), (25576,-0.791412), (25577,-0.973901), (25578,-1.030974), (25579,-0.810750), (25580,-0.802332), (25581,-0.975065), (25582,-1.026102), (25583,-1.179793), (25584,-0.888962), (25585,-1.023612), (25586,-1.044918), (25587,-0.804719), (25588,-0.640236), (25589,-0.788348), (25590,-0.873298), (25591,-0.909470), (25592,-0.557324), (25593,-0.712875), (25594,-0.791320), (25595,-0.926426), (25596,-0.492998), (25597,-0.647616), (25598,-0.692617), (25599,-0.875569), (25600,-0.609358), (25601,-0.745398), (25602,-0.812696), (25603,-0.972887), (25604,-0.437268), (25605,-0.593746), (25606,-0.663831), (25607,-0.807766), (25608,-0.595438), (25609,-0.753769), (25610,-0.807129), (25611,-0.941315), (25612,-0.532501), (25613,-0.688979), (25614,-0.746522), (25615,-0.913219), (25616,-0.637252), (25617,-0.773292), (25618,-0.832688), (25619,-0.985916), (25620,-0.460047), (25621,-0.621640), (25622,-0.678250), (25623,-0.841697), (25624,-0.679994), (25625,-0.716166), (25626,-0.889832), (25627,-0.882804), (25628,-0.637495), (25629,-0.674600), (25630,-0.874741), (25631,-0.589482), (25632,-0.760825), (25633,-0.845306), (25634,-0.985991), (25635,-0.833117), (25636,-0.590595), (25637,-0.663460), (25638,-0.792067), (25639,-0.522143), (25640,-0.833760), (25641,-0.914528), (25642,-1.115595), (25643,-0.666374), (25644,-0.816809), (25645,-0.893394), (25646,-1.002033), (25647,-0.789704), (25648,-0.950821), (25649,-0.997219), (25650,-1.121179), (25651,-0.591133), (25652,-0.726709), (25653,-0.771710), (25654,-0.938870), (25655,-0.551891), (25656,-0.682821), (25657,-0.721779), (25658,-0.876404), (25659,-0.849402), (25660,-0.599446), (25661,-0.681141), (25662,-0.838088), (25663,-0.542147), (25664,-0.714417), (25665,-0.747802), (25666,-0.896384), (25667,-0.750009), (25668,-0.524212), (25669,-0.572462), (25670,-0.743805), (25671,-0.458547), (25672,-0.609915), (25673,-0.653056), (25674,-0.843441), (25675,-0.857784), (25676,-0.613866), (25677,-0.642148), (25678,-0.807911), (25679,-0.529622), (25680,-0.732549), (25681,-0.730174), (25682,-0.904303), (25683,-0.792299), (25684,-0.518193), (25685,-0.592918), (25686,-0.783772), (25687,-0.459497), (25688,-0.607146), (25689,-0.666548), (25690,-0.839745), (25691,-0.829004), (25692,-0.612029), (25693,-0.628696), (25694,-0.822331), (25695,-0.570059), (25696,-0.729323), (25697,-0.765031), (25698,-0.915936), (25699,-0.779317), (25700,-0.496845), (25701,-0.571107), (25702,-0.724798), (25703,-0.429790), (25704,-0.745126), (25705,-0.791517), (25706,-0.963787), (25707,-0.557760), (25708,-0.703091), (25709,-0.788505), (25710,-0.932904), (25711,-0.688522), (25712,-0.828744), (25713,-0.876062), (25714,-1.070166), (25715,-0.513645), (25716,-0.648295), (25717,-0.703508), (25718,-0.854413), (25719,-0.500877), (25720,-0.902606), (25721,-0.958289), (25722,-1.104084), (25723,-0.692021), (25724,-0.856394), (25725,-0.919510), (25726,-1.083420), (25727,-0.829746), (25728,-1.115821), (25729,-1.149207), (25730,-1.294539), (25731,-0.738945), (25732,-0.913074), (25733,-0.947393), (25734,-1.112693), (25735,-0.763804), (25736,-1.046623), (25737,-1.109732), (25738,-1.242992), (25739,-0.849507), (25740,-0.989723), (25741,-1.062594), (25742,-1.177269), (25743,-0.968190), (25744,-1.119558), (25745,-1.191497), (25746,-1.325676), (25747,-0.776589), (25748,-0.891263), (25749,-0.936264), (25750,-1.118753), (25751,-0.773113), (25752,-0.773055), (25753,-0.942075), (25754,-1.005191), (25755,-1.154236), (25756,-0.751928), (25757,-0.909795), (25758,-0.944114), (25759,-1.094549), (25760,-0.823692), (25761,-0.982030), (25762,-1.044213), (25763,-1.171893), (25764,-0.657645), (25765,-0.790898), (25766,-0.841466), (25767,-1.011882), (25768,-0.824631), (25769,-0.981108), (25770,-1.036792), (25771,-0.793343), (25772,-0.793285), (25773,-0.928397), (25774,-0.999409), (25775,-1.178648), (25776,-0.897103), (25777,-1.053117), (25778,-1.114373), (25779,-0.889966), (25780,-0.757530), (25781,-0.903325), (25782,-0.959472), (25783,-1.009582), (25784,-0.998372), (25785,-1.142777), (25786,-1.178022), (25787,-0.938286), (25788,-0.888060), (25789,-1.051970), (25790,-1.123445), (25791,-1.285965), (25792,-1.007213), (25793,-1.156258), (25794,-1.191966), (25795,-0.945724), (25796,-0.798423), (25797,-1.009246), (25798,-1.051924), (25799,-1.125722), (25800,-0.873444), (25801,-1.022025), (25802,-1.101397), (25803,-0.848192), (25804,-0.821196), (25805,-1.000898), (25806,-1.038003), (25807,-1.227455), (25808,-0.925014), (25809,-1.094034), (25810,-1.162723), (25811,-0.949461), (25812,-0.790087), (25813,-0.968856), (25814,-1.038478), (25815,-1.092765), (25816,-0.820049), (25817,-0.964917), (25818,-1.021528), (25819,-1.192401), (25820,-0.802635), (25821,-0.945180), (25822,-0.979493), (25823,-1.102063), (25824,-0.840036), (25825,-0.972356), (25826,-1.032685), (25827,-1.172907), (25828,-0.621490), (25829,-0.796552), (25830,-0.877783), (25831,-1.019396), (25832,-0.679792), (25833,-0.854848), (25834,-0.881271), (25835,-1.054467), (25836,-0.639617), (25837,-0.784949), (25838,-0.804402), (25839,-0.973422), (25840,-0.720211), (25841,-0.865079), (25842,-0.930981), (25843,-1.065625), (25844,-0.509104), (25845,-0.658149), (25846,-0.727771), (25847,-0.907010), (25848,-0.580875), (25849,-0.707159), (25850,-0.759129), (25851,-0.952763), (25852,-0.542560), (25853,-0.678599), (25854,-0.738465), (25855,-0.903302), (25856,-0.619903), (25857,-0.748974), (25858,-0.816272), (25859,-0.958348), (25860,-0.406011), (25861,-0.553659), (25862,-0.620488), (25863,-0.792764), (25864,-0.608300), (25865,-0.732730), (25866,-0.791200), (25867,-0.950927), (25868,-0.543046), (25869,-0.705097), (25870,-0.765890), (25871,-0.920971), (25872,-0.690527), (25873,-0.803342), (25874,-0.860416), (25875,-1.000175), (25876,-0.462233), (25877,-0.612204), (25878,-0.684613), (25879,-0.844340), (25880,-0.680320), (25881,-0.736467), (25882,-0.871573), (25883,-0.917037), (25884,-0.657796), (25885,-0.707437), (25886,-0.863915), (25887,-0.603741), (25888,-0.795985), (25889,-0.846559), (25890,-0.990494), (25891,-0.852022), (25892,-0.606713), (25893,-0.697230), (25894,-0.825837), (25895,-0.535938), (25896,-0.740255), (25897,-0.818700), (25898,-0.970068), (25899,-0.929603), (25900,-0.686611), (25901,-0.767842), (25902,-0.866725), (25903,-0.582863), (25904,-0.750023), (25905,-0.801060), (25906,-0.972403), (25907,-0.817205), (25908,-0.571427), (25909,-0.649408), (25910,-0.857444), (25911,-0.526670), (25912,-0.706835), (25913,-0.752763), (25914,-0.886016), (25915,-0.873879), (25916,-0.634143), (25917,-0.676821), (25918,-0.839804), (25919,-0.561052), (25920,-0.759332), (25921,-0.782499), (25922,-0.972420), (25923,-0.818619), (25924,-0.552402), (25925,-0.635493), (25926,-0.814732), (25927,-0.524364), (25928,-0.684561), (25929,-0.750927), (25930,-0.916227), (25931,-0.865080), (25932,-0.614192), (25933,-0.663839), (25934,-0.853297), (25935,-0.564788), (25936,-0.747277), (25937,-0.777876), (25938,-0.936677), (25939,-0.777297), (25940,-0.522232), (25941,-0.602067), (25942,-0.769696), (25943,-0.486761), (25944,-0.674359), (25945,-0.711927), (25946,-0.856326), (25947,-0.850232), (25948,-0.616538), (25949,-0.653174), (25950,-0.837985), (25951,-0.545764), (25952,-0.726393), (25953,-0.760711), (25954,-0.936694), (25955,-0.778247), (25956,-0.522256), (25957,-0.572829), (25958,-0.748812), (25959,-0.472846), (25960,-0.705040), (25961,-0.777442), (25962,-0.979442), (25963,-0.589670), (25964,-0.749403), (25965,-0.765600), (25966,-0.908609), (25967,-0.659117), (25968,-0.805846), (25969,-0.875925), (25970,-1.005928), (25971,-0.443828), (25972,-0.642115), (25973,-0.696865), (25974,-0.833838), (25975,-0.481692), (25976,-0.912224), (25977,-0.973011), (25978,-1.129495), (25979,-0.737400), (25980,-0.889701), (25981,-0.941201), (25982,-1.105111), (25983,-0.836578), (25984,-1.054833), (25985,-1.094725), (25986,-1.233551), (25987,-0.714650), (25988,-0.881347), (25989,-0.918915), (25990,-1.060064), (25991,-0.709315), (25992,-0.877408), (25993,-1.027843), (25994,-1.061228), (25995,-0.841467), (25996,-0.832586), (25997,-1.009965), (25998,-1.020126), (25999,-1.223523), (26000,-0.996329), (26001,-1.151873), (26002,-1.231245), (26003,-0.969680), (26004,-0.807051), (26005,-0.949590), (26006,-0.989018), (26007,-1.075822), (26008,-0.904369), (26009,-1.033439), (26010,-1.072861), (26011,-0.831272), (26012,-0.784765), (26013,-0.964930), (26014,-1.008535), (26015,-1.193816), (26016,-0.923423), (26017,-1.082223), (26018,-1.114212), (26019,-0.898634), (26020,-0.755509), (26021,-0.905024), (26022,-0.972316), (26023,-1.028000), (26024,-0.785014), (26025,-0.939632), (26026,-0.980450), (26027,-0.755116), (26028,-0.775959), (26029,-0.885524), (26030,-0.942598), (26031,-1.119977), (26032,-0.839364), (26033,-1.005598), (26034,-1.085902), (26035,-0.826191), (26036,-0.679817), (26037,-0.827935), (26038,-0.840882), (26039,-0.961599), (26040,-0.944353), (26041,-1.077143), (26042,-1.143972), (26043,-0.887981), (26044,-0.880490), (26045,-1.049510), (26046,-1.108443), (26047,-1.271890), (26048,-0.988028), (26049,-1.098056), (26050,-1.163489), (26051,-0.960452), (26052,-0.762983), (26053,-0.931076), (26054,-0.973284), (26055,-1.063807), (26056,-0.804560), (26057,-0.967543), (26058,-1.017184), (26059,-0.768625), (26060,-0.752775), (26061,-0.907856), (26062,-0.970509), (26063,-1.159034), (26064,-0.858453), (26065,-1.011211), (26066,-1.054822), (26067,-0.824835), (26068,-0.676144), (26069,-0.859559), (26070,-0.880873), (26071,-0.927727), (26072,-0.827808), (26073,-1.018656), (26074,-1.013488), (26075,-0.788154), (26076,-0.751402), (26077,-0.936214), (26078,-0.992824), (26079,-1.198074), (26080,-0.872409), (26081,-1.036782), (26082,-1.132409), (26083,-0.863876), (26084,-0.723544), (26085,-0.853547), (26086,-0.964965), (26087,-1.028545), (26088,-0.734927), (26089,-0.858887), (26090,-0.929436), (26091,-0.654866), (26092,-0.636693), (26093,-0.804317), (26094,-0.898090), (26095,-1.051781), (26096,-0.750267), (26097,-0.908135), (26098,-0.964282), (26099,-0.718046), (26100,-0.578641), (26101,-0.765775), (26102,-0.819599), (26103,-0.891538), (26104,-0.500376), (26105,-0.643384), (26106,-0.694885), (26107,-0.860655), (26108,-0.478785), (26109,-0.624580), (26110,-0.676081), (26111,-0.848350), (26112,-0.608151), (26113,-0.711673), (26114,-0.754351), (26115,-0.921511), (26116,-0.369174), (26117,-0.502890), (26118,-0.632893), (26119,-0.768469), (26120,-0.562640), (26121,-0.700539), (26122,-0.748327), (26123,-0.895975), (26124,-0.534080), (26125,-0.677552), (26126,-0.717907), (26127,-0.845118), (26128,-0.577517), (26129,-0.733062), (26130,-0.804074), (26131,-0.966124), (26132,-0.396598), (26133,-0.580483), (26134,-0.635233), (26135,-0.764310), (26136,-0.631404), (26137,-0.695917), (26138,-0.848211), (26139,-0.806350), (26140,-0.564291), (26141,-0.609756), (26142,-0.782025), (26143,-0.493517), (26144,-0.684834), (26145,-0.731225), (26146,-0.896062), (26147,-0.739005), (26148,-0.497416), (26149,-0.532191), (26150,-0.704467), (26151,-0.441507), (26152,-0.801432), (26153,-0.839464), (26154,-1.001051), (26155,-0.595957), (26156,-0.717131), (26157,-0.817867), (26158,-0.942761), (26159,-0.681660), (26160,-0.845570), (26161,-0.914722), (26162,-1.062371), (26163,-0.510497), (26164,-0.639567), (26165,-0.718011), (26166,-0.891214), (26167,-0.521417), (26168,-0.634695), (26169,-0.682946), (26170,-0.877050), (26171,-0.856553), (26172,-0.638652), (26173,-0.676220), (26174,-0.802967), (26175,-0.496344), (26176,-0.665364), (26177,-0.733589), (26178,-0.932803), (26179,-0.768777), (26180,-0.558771), (26181,-0.605625), (26182,-0.736555), (26183,-0.450370), (26184,-0.648187), (26185,-0.662994), (26186,-0.813899), (26187,-0.841248), (26188,-0.578288), (26189,-0.634435), (26190,-0.812740), (26191,-0.544670), (26192,-0.715086), (26193,-0.749868), (26194,-0.886371), (26195,-0.734424), (26196,-0.497474), (26197,-0.570809), (26198,-0.711958), (26199,-0.438778), (26200,-0.613371), (26201,-0.663945), (26202,-0.809276), (26203,-0.787384), (26204,-0.527679), (26205,-0.619123), (26206,-0.799295), (26207,-0.494062), (26208,-0.667264), (26209,-0.689504), (26210,-0.873383), (26211,-0.732587), (26212,-0.463121), (26213,-0.514628), (26214,-0.705476), (26215,-0.427650), (26216,-0.620357), (26217,-0.743861), (26218,-0.787929), (26219,-0.531468), (26220,-0.510045), (26221,-0.676278), (26222,-0.723139), (26223,-0.913523), (26224,-0.636624), (26225,-0.820046), (26226,-0.853431), (26227,-0.614159), (26228,-0.458962), (26229,-0.592215), (26230,-0.642788), (26231,-0.695685), (26232,-0.791312), (26233,-0.856751), (26234,-1.034593), (26235,-0.622530), (26236,-0.773434), (26237,-0.833301), (26238,-1.006960), (26239,-0.804851), (26240,-0.991985), (26241,-1.154969), (26242,-1.231554), (26243,-0.981129), (26244,-0.775306), (26245,-0.935497), (26246,-1.005112), (26247,-1.043144), (26248,-0.869368), (26249,-1.004481), (26250,-1.076420), (26251,-0.832501), (26252,-0.810615), (26253,-0.979171), (26254,-1.000948), (26255,-1.212697), (26256,-0.931621), (26257,-1.077416), (26258,-1.093150), (26259,-0.875712), (26260,-0.745129), (26261,-0.890461), (26262,-0.937785), (26263,-1.037131), (26264,-0.751410), (26265,-0.882803), (26266,-0.928731), (26267,-1.086135), (26268,-0.705198), (26269,-0.849133), (26270,-0.927572), (26271,-1.094738), (26272,-0.814589), (26273,-0.949702), (26274,-1.009562), (26275,-1.154430), (26276,-0.629957), (26277,-0.763210), (26278,-0.814247), (26279,-0.974444), (26280,-0.779761), (26281,-0.882357), (26282,-0.956618), (26283,-0.718742), (26284,-0.690350), (26285,-0.847297), (26286,-0.905761), (26287,-1.090109), (26288,-0.781632), (26289,-0.966444), (26290,-1.028627), (26291,-0.787501), (26292,-0.626724), (26293,-0.787385), (26294,-0.829130), (26295,-0.903861), (26296,-0.902407), (26297,-1.050525), (26298,-1.105282), (26299,-0.861826), (26300,-0.828794), (26301,-1.011283), (26302,-1.044205), (26303,-1.210438), (26304,-0.927966), (26305,-1.092340), (26306,-1.143377), (26307,-0.891099), (26308,-0.755876), (26309,-0.898421), (26310,-0.966641), (26311,-1.057164), (26312,-0.792807), (26313,-0.943712), (26314,-0.986390), (26315,-0.735038), (26316,-0.724298), (26317,-0.884495), (26318,-0.947147), (26319,-1.124063), (26320,-0.813257), (26321,-0.994355), (26322,-1.055142), (26323,-0.807047), (26324,-0.629552), (26325,-0.797181), (26326,-0.861224), (26327,-0.889963), (26328,-0.653483), (26329,-0.828539), (26330,-0.868894), (26331,-1.036054), (26332,-0.666257), (26333,-0.802296), (26334,-0.871918), (26335,-1.018640), (26336,-0.766825), (26337,-0.886146), (26338,-0.932537), (26339,-1.114562), (26340,-0.539927), (26341,-0.693618), (26342,-0.790177), (26343,-0.908565), (26344,-0.893642), (26345,-0.603744), (26346,-0.769977), (26347,-0.847952), (26348,-0.583138), (26349,-0.578434), (26350,-0.734448), (26351,-0.796167), (26352,-0.967047), (26353,-0.665533), (26354,-0.811328), (26355,-0.874901), (26356,-0.613800), (26357,-0.433982), (26358,-0.615081), (26359,-0.697702), (26360,-0.493269), (26361,-0.643710), (26362,-0.681742), (26363,-0.839146), (26364,-0.431266), (26365,-0.587743), (26366,-0.658292), (26367,-0.801764), (26368,-0.601971), (26369,-0.757058), (26370,-0.806236), (26371,-0.934843), (26372,-0.400620), (26373,-0.570103), (26374,-0.613708), (26375,-0.767862), (26376,-0.889043), (26377,-0.616327), (26378,-0.768621), (26379,-0.835450), (26380,-0.585495), (26381,-0.580334), (26382,-0.737738), (26383,-0.790172), (26384,-0.954545), (26385,-0.673933), (26386,-0.840166), (26387,-0.899563), (26388,-0.644498), (26389,-0.470723), (26390,-0.636956), (26391,-0.675451), (26392,-0.740421), (26393,-0.781702), (26394,-0.899163), (26395,-0.935805), (26396,-0.683990), (26397,-0.736887), (26398,-0.905907), (26399,-0.624368), (26400,-0.793387), (26401,-0.877868), (26402,-1.032023), (26403,-0.873106), (26404,-0.624084), (26405,-0.707632), (26406,-0.855750), (26407,-0.576071), (26408,-0.595518), (26409,-0.744569), (26410,-0.779344), (26411,-0.950224), (26412,-0.537234), (26413,-0.683490), (26414,-0.749391), (26415,-0.881251), (26416,-0.615504), (26417,-0.769659), (26418,-0.824877), (26419,-1.021301), (26420,-0.463851), (26421,-0.623116), (26422,-0.679263), (26423,-0.799510), (26424,-0.633164), (26425,-0.691634), (26426,-0.859259), (26427,-0.812754), (26428,-0.593920), (26429,-0.662143), (26430,-0.830698), (26431,-0.523146), (26432,-0.696810), (26433,-0.770608), (26434,-0.907113), (26435,-0.766778), (26436,-0.554912), (26437,-0.612917), (26438,-0.758711), (26439,-0.508292), (26440,-0.586270), (26441,-0.728814), (26442,-0.777064), (26443,-0.910318), (26444,-0.514511), (26445,-0.677957), (26446,-0.729923), (26447,-0.884543), (26448,-0.613686), (26449,-0.780847), (26450,-0.842104), (26451,-1.000439), (26452,-0.477362), (26453,-0.581816), (26454,-0.634712), (26455,-0.786081), (26456,-0.693124), (26457,-0.761813), (26458,-0.906214), (26459,-0.921486), (26460,-0.676640), (26461,-0.730000), (26462,-0.909239), (26463,-0.621660), (26464,-0.753519), (26465,-0.786442), (26466,-0.975899), (26467,-0.852751), (26468,-0.613479), (26469,-0.672878), (26470,-0.860012), (26471,-0.562214), (26472,-0.606749), (26473,-0.749292), (26474,-0.806368), (26475,-0.591714), (26476,-0.533132), (26477,-0.718408), (26478,-0.778271), (26479,-0.990953), (26480,-0.715915), (26481,-0.863568), (26482,-0.895097), (26483,-0.638174), (26484,-0.489015), (26485,-0.643635), (26486,-0.679344), (26487,-0.767076), (26488,-0.726609), (26489,-0.893770), (26490,-0.962923), (26491,-0.752915), (26492,-0.743568), (26493,-0.908407), (26494,-0.944581), (26495,-1.136824), (26496,-0.860858), (26497,-0.984357), (26498,-1.028427), (26499,-1.155177), (26500,-0.579147), (26501,-0.750489), (26502,-0.815461), (26503,-0.944069), (26504,-0.838108), (26505,-0.969503), (26506,-1.012179), (26507,-0.786843), (26508,-0.797005), (26509,-0.956734), (26510,-1.005450), (26511,-1.171218), (26512,-0.891535), (26513,-1.087030), (26514,-1.127849), (26515,-0.869069), (26516,-0.705974), (26517,-0.838763), (26518,-0.910238), (26519,-0.990539), (26520,-0.669981), (26521,-0.839000), (26522,-0.869600), (26523,-0.999602), (26524,-0.617266), (26525,-0.780247), (26526,-0.868444), (26527,-1.000304), (26528,-0.772644), (26529,-0.896143), (26530,-0.958793), (26531,-1.147786), (26532,-0.651185), (26533,-0.793727), (26534,-0.854519), (26535,-1.017035), (26536,-0.892494), (26537,-1.066623), (26538,-1.105119), (26539,-0.857952), (26540,-0.852785), (26541,-0.988825), (26542,-1.036147), (26543,-1.226068), (26544,-0.939418), (26545,-1.073136), (26546,-1.121387), (26547,-0.903017), (26548,-0.762219), (26549,-0.908013), (26550,-0.936755), (26551,-0.981754), (26552,-0.761992), (26553,-0.885026), (26554,-0.931883), (26555,-1.077678), (26556,-0.663292), (26557,-0.834169), (26558,-0.932120), (26559,-1.076521), (26560,-0.809380), (26561,-0.953781), (26562,-0.989490), (26563,-1.140859), (26564,-0.616388), (26565,-0.790981), (26566,-0.814613), (26567,-0.984562), (26568,-0.801029), (26569,-0.992809), (26570,-1.076361), (26571,-0.849631), (26572,-0.823098), (26573,-0.981898), (26574,-1.027362), (26575,-1.186162), (26576,-0.899977), (26577,-1.075964), (26578,-1.136291), (26579,-0.895626), (26580,-0.733461), (26581,-0.855566), (26582,-0.903816), (26583,-0.980866), (26584,-0.715118), (26585,-0.874847), (26586,-0.910557), (26587,-1.084221), (26588,-0.670299), (26589,-0.820275), (26590,-0.909400), (26591,-1.009674), (26592,-0.738353), (26593,-0.887863), (26594,-0.940759), (26595,-1.112565), (26596,-0.592739), (26597,-0.745501), (26598,-0.812331), (26599,-0.940475), (26600,-0.914871), (26601,-0.629150), (26602,-0.773551), (26603,-0.846885), (26604,-0.625264), (26605,-0.601518), (26606,-0.783078), (26607,-0.789524), (26608,-0.991988), (26609,-0.708589), (26610,-0.827443), (26611,-0.932826), (26612,-0.678691), (26613,-0.509094), (26614,-0.683687), (26615,-0.717538), (26616,-0.619938), (26617,-0.759693), (26618,-0.813518), (26619,-0.979286), (26620,-0.574654), (26621,-0.730203), (26622,-0.778454), (26623,-0.949331), (26624,-1.341307), (26625,-1.084385), (26626,-1.208813), (26627,-0.857134), (26628,-0.988529), (26629,-0.878387), (26630,-1.055303), (26631,-1.010654), (26632,-1.326918), (26633,-1.052346), (26634,-1.169805), (26635,-0.839958), (26636,-0.981572), (26637,-1.016352), (26638,-1.195126), (26639,-1.274962), (26640,-1.430046), (26641,-1.145719), (26642,-1.304983), (26643,-0.961201), (26644,-1.108853), (26645,-0.955049), (26646,-1.088302), (26647,-1.068737), (26648,-0.869876), (26649,-1.032857), (26650,-1.081572), (26651,-1.252913), (26652,-0.842708), (26653,-0.968994), (26654,-1.010277), (26655,-1.180690), (26656,-0.942347), (26657,-1.036583), (26658,-1.099233), (26659,-1.247814), (26660,-0.682003), (26661,-0.849629), (26662,-0.902060), (26663,-1.052964), (26664,-0.972550), (26665,-1.145284), (26666,-1.191677), (26667,-0.977488), (26668,-0.959781), (26669,-1.114866), (26670,-1.171942), (26671,-1.327026), (26672,-1.045021), (26673,-1.222865), (26674,-1.279477), (26675,-1.019303), (26676,-0.843668), (26677,-1.005719), (26678,-1.053041), (26679,-1.139845), (26680,-0.969318), (26681,-1.111861), (26682,-1.127598), (26683,-0.904119), (26684,-0.911029), (26685,-1.088410), (26686,-1.136196), (26687,-1.300105), (26688,-1.033893), (26689,-1.177365), (26690,-1.214004), (26691,-0.987738), (26692,-0.823715), (26693,-0.996914), (26694,-1.027514), (26695,-1.097596), (26696,-0.924283), (26697,-1.112346), (26698,-1.179177), (26699,-0.947802), (26700,-0.907334), (26701,-1.055915), (26702,-1.109740), (26703,-1.303377), (26704,-1.015334), (26705,-1.141619), (26706,-1.160142), (26707,-0.924123), (26708,-0.816303), (26709,-0.987180), (26710,-1.015457), (26711,-1.113873), (26712,-0.793315), (26713,-0.939575), (26714,-0.998044), (26715,-1.145232), (26716,-0.715054), (26717,-0.865028), (26718,-0.924427), (26719,-1.073937), (26720,-0.834666), (26721,-0.982318), (26722,-1.080270), (26723,-1.246037), (26724,-0.691839), (26725,-0.832988), (26726,-0.868698), (26727,-1.012634), (26728,-0.850004), (26729,-1.025062), (26730,-1.070061), (26731,-0.795488), (26732,-0.807043), (26733,-0.941690), (26734,-1.005269), (26735,-1.154779), (26736,-0.886709), (26737,-1.035755), (26738,-1.103515), (26739,-0.846592), (26740,-0.720658), (26741,-0.903147), (26742,-0.952327), (26743,-1.041453), (26744,-0.977761), (26745,-1.111014), (26746,-1.147187), (26747,-0.919064), (26748,-0.888815), (26749,-1.062479), (26750,-1.134419), (26751,-1.291361), (26752,-1.623882), (26753,-1.355348), (26754,-1.136979), (26755,-1.158753), (26756,-1.322663), (26757,-1.126590), (26758,-1.198065), (26759,-1.256534), (26760,-1.517059), (26761,-1.235983), (26762,-0.979061), (26763,-1.044033), (26764,-1.194937), (26765,-1.201848), (26766,-1.377834), (26767,-1.451167), (26768,-1.620651), (26769,-1.330286), (26770,-1.072434), (26771,-1.134619), (26772,-1.277627), (26773,-1.111281), (26774,-1.212949), (26775,-1.242620), (26776,-1.537053), (26777,-1.250402), (26778,-1.013918), (26779,-1.070530), (26780,-1.194028), (26781,-1.196759), (26782,-1.357417), (26783,-1.401487), (26784,-1.558894), (26785,-1.266205), (26786,-1.038082), (26787,-1.062643), (26788,-1.205187), (26789,-1.064852), (26790,-1.147011), (26791,-1.198048), (26792,-1.389363), (26793,-1.091566), (26794,-0.823960), (26795,-0.881036), (26796,-1.070028), (26797,-1.056037), (26798,-1.236204), (26799,-1.284455), (26800,-1.478556), (26801,-1.214202), (26802,-0.932198), (26803,-0.967442), (26804,-1.141571), (26805,-0.987766), (26806,-1.069925), (26807,-1.106099), (26808,-1.534770), (26809,-1.259733), (26810,-1.010242), (26811,-1.056635), (26812,-1.227513), (26813,-1.243249), (26814,-1.425738), (26815,-1.430791), (26816,-1.569618), (26817,-1.311767), (26818,-1.045090), (26819,-1.084980), (26820,-1.232168), (26821,-1.138747), (26822,-1.190249), (26823,-1.260331), (26824,-1.414951), (26825,-1.134340), (26826,-0.883456), (26827,-0.934494), (26828,-1.118377), (26829,-1.089057), (26830,-1.284088), (26831,-1.353241), (26832,-1.506467), (26833,-1.249080), (26834,-0.978687), (26835,-1.028796), (26836,-1.181093), (26837,-1.003600), (26838,-1.059747), (26839,-1.125184), (26840,-1.496723), (26841,-1.201247), (26842,-0.960582), (26843,-1.024626), (26844,-1.177852), (26845,-1.167576), (26846,-1.353782), (26847,-1.372769), (26848,-1.536679), (26849,-1.261642), (26850,-0.988927), (26851,-1.051112), (26852,-1.228957), (26853,-1.080726), (26854,-1.161956), (26855,-1.206490), (26856,-1.283540), (26857,-1.420045), (26858,-0.748328), (26859,-0.904342), (26860,-0.967457), (26861,-1.118361), (26862,-1.109013), (26863,-1.260382), (26864,-1.314207), (26865,-1.460465), (26866,-0.785498), (26867,-0.945228), (26868,-1.020419), (26869,-1.165284), (26870,-0.940412), (26871,-1.099213), (26872,-1.199022), (26873,-0.954176), (26874,-1.099042), (26875,-0.739931), (26876,-0.867146), (26877,-0.881953), (26878,-1.033786), (26879,-1.123376), (26880,-1.256629), (26881,-0.945826), (26882,-1.116239), (26883,-0.760379), (26884,-0.909425), (26885,-0.778381), (26886,-0.942290), (26887,-0.905539), (26888,-1.107537), (26889,-1.272840), (26890,-0.987119), (26891,-0.722301), (26892,-0.786809), (26893,-0.957685), (26894,-0.936727), (26895,-1.110391), (26896,-1.178150), (26897,-1.333235), (26898,-1.038224), (26899,-0.817068), (26900,-0.852777), (26901,-1.019938), (26902,-0.859166), (26903,-0.929248), (26904,-0.851156), (26905,-1.024821), (26906,-1.056349), (26907,-0.827297), (26908,-0.850464), (26909,-1.038064), (26910,-1.098391), (26911,-1.265088), (26912,-0.964968), (26913,-1.136309), (26914,-1.193850), (26915,-0.940644), (26916,-0.748286), (26917,-0.925666), (26918,-0.972988), (26919,-1.006839), (26920,-1.339360), (26921,-1.061071), (26922,-0.838057), (26923,-0.898385), (26924,-1.028387), (26925,-0.992099), (26926,-1.184807), (26927,-1.246993), (26928,-1.394645), (26929,-1.139117), (26930,-0.912387), (26931,-0.971785), (26932,-1.112005), (26933,-0.972600), (26934,-1.061262), (26935,-1.089075), (26936,-0.863274), (26937,-1.077813), (26938,-1.113987), (26939,-0.862174), (26940,-0.858402), (26941,-1.016273), (26942,-1.071491), (26943,-1.252587), (26944,-0.966402), (26945,-1.112196), (26946,-1.163234), (26947,-0.887267), (26948,-0.765513), (26949,-0.903411), (26950,-0.964667), (26951,-1.017098), (26952,-1.156390), (26953,-0.893894), (26954,-1.058268), (26955,-0.746535), (26956,-0.890007), (26957,-0.868119), (26958,-1.025991), (26959,-1.103969), (26960,-1.232113), (26961,-0.987732), (26962,-1.142352), (26963,-0.792995), (26964,-0.896056), (26965,-0.771979), (26966,-0.942392), (26967,-0.912143), (26968,-0.815472), (26969,-0.960802), (26970,-1.028561), (26971,-0.758633), (26972,-0.753931), (26973,-0.897868), (26974,-0.954479), (26975,-1.138827), (26976,-0.848461), (26977,-1.009584), (26978,-1.042506), (26979,-0.816240), (26980,-0.667081), (26981,-0.834707), (26982,-0.880170), (26983,-0.962329), (26984,-1.233537), (26985,-0.944564), (26986,-0.677888), (26987,-0.758653), (26988,-0.903054), (26989,-0.930867), (26990,-1.091525), (26991,-1.174613), (26992,-1.330627), (26993,-1.028648), (26994,-0.790305), (26995,-0.837627), (26996,-0.994105), (26997,-0.859345), (26998,-0.919208), (26999,-0.988825), (27000,-1.413316), (27001,-1.115983), (27002,-0.858132), (27003,-0.907312), (27004,-1.064718), (27005,-1.084171), (27006,-1.257370), (27007,-1.317233), (27008,-1.269798), (27009,-1.410947), (27010,-1.059732), (27011,-1.195308), (27012,-1.021530), (27013,-1.187763), (27014,-1.168662), (27015,-1.359977), (27016,-1.485333), (27017,-1.200077), (27018,-0.935258), (27019,-0.995586), (27020,-1.172966), (27021,-1.137607), (27022,-1.309878), (27023,-1.336298), (27024,-1.494634), (27025,-1.206590), (27026,-0.980324), (27027,-1.044368), (27028,-1.210600), (27029,-1.088846), (27030,-1.138954), (27031,-1.194173), (27032,-1.332070), (27033,-1.077006), (27034,-1.232555), (27035,-0.896204), (27036,-1.063365), (27037,-1.053090), (27038,-1.212355), (27039,-1.299158), (27040,-1.436592), (27041,-1.174095), (27042,-1.336148), (27043,-0.991436), (27044,-1.133514), (27045,-0.952305), (27046,-1.093919), (27047,-1.098042), (27048,-1.406410), (27049,-1.122547), (27050,-0.899068), (27051,-0.938029), (27052,-1.057347), (27053,-1.050788), (27054,-1.235135), (27055,-1.296856), (27056,-1.463553), (27057,-1.150427), (27058,-0.890718), (27059,-0.921317), (27060,-1.131212), (27061,-0.970905), (27062,-1.018691), (27063,-1.089237), (27064,-1.500258), (27065,-1.229401), (27066,-0.981304), (27067,-1.021658), (27068,-1.198574), (27069,-1.195730), (27070,-1.362891), (27071,-1.420896), (27072,-1.562975), (27073,-1.324632), (27074,-1.070962), (27075,-1.157301), (27076,-1.304489), (27077,-1.153007), (27078,-1.219837), (27079,-1.265301), (27080,-1.435713), (27081,-1.176005), (27082,-0.920940), (27083,-0.980803), (27084,-1.127991), (27085,-1.107961), (27086,-1.308101), (27087,-1.358210), (27088,-1.513759), (27089,-1.229431), (27090,-1.018494), (27091,-1.072783), (27092,-1.233441), (27093,-1.075457), (27094,-1.165512), (27095,-1.198434), (27096,-1.399039), (27097,-1.104957), (27098,-1.240533), (27099,-0.919510), (27100,-1.065769), (27101,-1.040630), (27102,-1.206862), (27103,-1.272763), (27104,-1.422738), (27105,-1.163493), (27106,-1.320436), (27107,-0.954357), (27108,-1.098758), (27109,-1.006731), (27110,-1.109792), (27111,-1.073505), (27112,-1.252279), (27113,-0.987460), (27114,-1.144403), (27115,-0.802942), (27116,-0.945949), (27117,-0.946357), (27118,-1.070321), (27119,-1.145512), (27120,-1.279694), (27121,-1.041352), (27122,-1.191791), (27123,-0.855904), (27124,-1.031891), (27125,-0.880409), (27126,-1.022023), (27127,-0.979233), (27128,-1.157078), (27129,-0.897369), (27130,-1.048273), (27131,-0.713315), (27132,-0.859110), (27133,-0.833505), (27134,-0.967223), (27135,-1.097690), (27136,-1.226762), (27137,-0.961943), (27138,-1.126317), (27139,-0.769993), (27140,-0.913001), (27141,-0.780563), (27142,-0.946331), (27143,-0.914224), (27144,-1.202154), (27145,-0.932226), (27146,-1.095671), (27147,-0.750030), (27148,-0.928339), (27149,-0.934321), (27150,-1.089870), (27151,-1.160881), (27152,-1.280664), (27153,-1.010736), (27154,-1.171394), (27155,-0.852229), (27156,-0.968296), (27157,-0.811240), (27158,-0.982117), (27159,-0.948152), (27160,-0.887247), (27161,-1.050228), (27162,-1.105910), (27163,-0.857349), (27164,-0.822919), (27165,-0.989152), (27166,-1.031364), (27167,-1.200848), (27168,-0.911875), (27169,-1.082288), (27170,-1.157015), (27171,-0.896841), (27172,-0.711451), (27173,-0.874432), (27174,-0.924076), (27175,-1.009022), (27176,-0.855682), (27177,-0.997296), (27178,-1.078061), (27179,-0.832286), (27180,-0.800644), (27181,-0.976631), (27182,-1.041139), (27183,-1.227344), (27184,-0.930475), (27185,-1.066515), (27186,-1.112908), (27187,-0.878746), (27188,-0.737947), (27189,-0.886994), (27190,-0.926883), (27191,-1.014151), (27192,-0.841767), (27193,-1.012180), (27194,-1.077152), (27195,-0.816979), (27196,-0.802058), (27197,-0.972935), (27198,-1.027688), (27199,-1.216216), (27200,-0.903090), (27201,-1.072110), (27202,-1.105497), (27203,-0.870406), (27204,-0.741219), (27205,-0.866111), (27206,-0.900892), (27207,-0.979799), (27208,-0.787906), (27209,-0.969931), (27210,-1.025149), (27211,-0.797026), (27212,-0.772815), (27213,-0.923254), (27214,-0.990550), (27215,-1.144240), (27216,-0.872454), (27217,-1.057730), (27218,-1.112949), (27219,-0.842091), (27220,-0.692932), (27221,-0.851732), (27222,-0.896731), (27223,-0.997005), (27224,-0.797216), (27225,-0.932792), (27226,-0.995442), (27227,-0.760815), (27228,-0.762616), (27229,-0.900979), (27230,-0.949230), (27231,-1.128468), (27232,-0.860862), (27233,-0.995973), (27234,-1.036327), (27235,-0.794733), (27236,-0.643716), (27237,-0.831315), (27238,-0.842871), (27239,-0.923636), (27240,-0.840899), (27241,-0.989945), (27242,-0.660562), (27243,-0.794743), (27244,-0.792829), (27245,-0.934443), (27246,-1.017531), (27247,-1.170757), (27248,-0.903151), (27249,-1.042907), (27250,-0.738142), (27251,-0.922025), (27252,-0.764504), (27253,-0.920053), (27254,-0.901882), (27255,-1.061146), (27256,-1.041117), (27257,-1.190162), (27258,-0.861244), (27259,-0.980097), (27260,-0.947062), (27261,-1.101681), (27262,-1.196846), (27263,-1.362149), (27264,-1.449417), (27265,-1.178560), (27266,-0.926747), (27267,-0.988468), (27268,-1.158417), (27269,-0.993464), (27270,-1.085842), (27271,-1.157782), (27272,-1.374179), (27273,-1.106109), (27274,-0.874270), (27275,-0.945280), (27276,-1.067386), (27277,-1.035278), (27278,-1.197331), (27279,-1.282276), (27280,-1.435038), (27281,-1.155356), (27282,-0.946276), (27283,-0.940646), (27284,-1.104091), (27285,-0.962828), (27286,-1.069604), (27287,-1.110888), (27288,-1.344008), (27289,-1.493518), (27290,-0.832020), (27291,-0.968990), (27292,-1.062296), (27293,-1.210878), (27294,-1.211286), (27295,-1.375195), (27296,-1.441561), (27297,-1.578066), (27298,-0.907279), (27299,-1.069331), (27300,-1.110614), (27301,-1.278704), (27302,-1.034323), (27303,-1.217742), (27304,-1.423456), (27305,-1.183256), (27306,-0.893819), (27307,-1.073986), (27308,-1.106908), (27309,-1.277321), (27310,-1.258220), (27311,-1.439316), (27312,-1.487567), (27313,-1.196736), (27314,-0.904512), (27315,-1.084215), (27316,-1.184489), (27317,-1.265719), (27318,-1.122598), (27319,-1.242380), (27320,-1.318965), (27321,-1.463366), (27322,-0.785612), (27323,-0.919330), (27324,-0.954574), (27325,-1.119878), (27326,-1.124466), (27327,-1.260971), (27328,-1.330587), (27329,-1.489388), (27330,-0.822781), (27331,-0.963931), (27332,-1.021936), (27333,-1.196994), (27334,-0.943323), (27335,-1.121167), (27336,-1.226551), (27337,-1.369558), (27338,-0.710849), (27339,-0.866398), (27340,-0.951343), (27341,-1.089706), (27342,-1.118448), (27343,-1.296756), (27344,-1.350581), (27345,-1.487086), (27346,-0.767063), (27347,-0.945372), (27348,-0.987119), (27349,-1.154745), (27350,-0.881565), (27351,-1.036186), (27352,-1.364526), (27353,-1.500102), (27354,-0.833031), (27355,-0.985793), (27356,-1.021038), (27357,-1.203527), (27358,-1.212760), (27359,-1.364129), (27360,-1.400767), (27361,-1.546562), (27362,-0.903180), (27363,-1.055942), (27364,-1.131133), (27365,-1.255561), (27366,-1.013967), (27367,-1.157903), (27368,-1.219624), (27369,-1.373315), (27370,-0.691381), (27371,-0.851110), (27372,-0.949061), (27373,-1.113900), (27374,-1.081793), (27375,-1.253135), (27376,-1.297670), (27377,-1.464366), (27378,-0.801940), (27379,-0.967708), (27380,-1.033610), (27381,-1.151534), (27382,-0.918766), (27383,-1.069205), (27384,-1.156473), (27385,-1.286475), (27386,-0.649596), (27387,-0.790281), (27388,-0.830635), (27389,-0.988971), (27390,-1.007959), (27391,-1.181158), (27392,-1.264246), (27393,-1.431872), (27394,-0.767588), (27395,-0.885977), (27396,-0.941195), (27397,-1.096279), (27398,-0.846325), (27399,-0.987475), (27400,-1.240103), (27401,-1.400296), (27402,-0.708607), (27403,-0.934295), (27404,-0.987655), (27405,-1.134843), (27406,-1.117600), (27407,-1.279187), (27408,-1.317683), (27409,-1.470445), (27410,-0.799194), (27411,-0.979825), (27412,-1.039688), (27413,-1.159007), (27414,-0.923451), (27415,-1.089684), (27416,-1.174164), (27417,-0.862896), (27418,-1.037954), (27419,-0.686275), (27420,-0.876661), (27421,-0.878462), (27422,-1.021934), (27423,-1.103628), (27424,-1.236417), (27425,-0.956270), (27426,-1.123431), (27427,-0.768965), (27428,-0.913366), (27429,-0.760955), (27430,-0.909072), (27431,-0.902512), (27432,-1.307959), (27433,-1.053824), (27434,-0.835920), (27435,-0.904608), (27436,-1.048080), (27437,-1.022476), (27438,-1.217507), (27439,-1.269938), (27440,-1.396224), (27441,-1.099355), (27442,-0.876805), (27443,-0.933416), (27444,-1.119622), (27445,-0.969069), (27446,-1.047512), (27447,-1.082292), (27448,-1.353035), (27449,-1.061741), (27450,-0.806677), (27451,-0.880010), (27452,-1.019766), (27453,-1.028999), (27454,-1.200805), (27455,-1.270422), (27456,-1.417146), (27457,-1.142573), (27458,-0.919559), (27459,-0.945049), (27460,-1.107565), (27461,-0.926356), (27462,-0.968103), (27463,-1.037256), (27464,-1.313574), (27465,-1.032033), (27466,-0.810413), (27467,-0.844264), (27468,-0.997491), (27469,-0.991860), (27470,-1.178994), (27471,-1.237464), (27472,-1.393477), (27473,-1.127730), (27474,-0.876381), (27475,-0.923238), (27476,-1.062995), (27477,-0.901758), (27478,-0.970446), (27479,-1.016375), (27480,-1.117577), (27481,-0.836502), (27482,-0.947923), (27483,-0.636190), (27484,-0.794062), (27485,-0.785644), (27486,-0.944444), (27487,-1.048899), (27488,-1.189584), (27489,-0.927552), (27490,-1.071489), (27491,-0.741177), (27492,-0.868391), (27493,-0.702045), (27494,-0.873387), (27495,-0.850106), (27496,-1.343807), (27497,-0.647473), (27498,-0.845290), (27499,-0.917695), (27500,-1.055128), (27501,-1.059252), (27502,-1.266825), (27503,-1.302534), (27504,-1.467837), (27505,-0.787296), (27506,-0.945631), (27507,-1.018036), (27508,-1.170333), (27509,-0.906908), (27510,-1.083359), (27511,-1.184097), (27512,-1.335466), (27513,-1.032559), (27514,-0.779817), (27515,-0.851292), (27516,-1.004054), (27517,-0.987740), (27518,-1.130747), (27519,-1.165992), (27520,-1.316896), (27521,-1.493347), (27522,-1.247108), (27523,-0.989257), (27524,-1.042618), (27525,-1.187483), (27526,-1.021601), (27527,-1.112121), (27528,-1.419095), (27529,-1.576967), (27530,-0.892709), (27531,-1.022711), (27532,-1.052382), (27533,-1.267851), (27534,-1.268722), (27535,-1.405692), (27536,-1.462303), (27537,-1.615530), (27538,-0.961000), (27539,-1.130949), (27540,-1.183380), (27541,-1.356579), (27542,-1.119630), (27543,-1.262173), (27544,-1.277445), (27545,-1.414414), (27546,-1.161672), (27547,-0.917755), (27548,-1.015242), (27549,-1.170791), (27550,-1.136362), (27551,-1.313742), (27552,-1.345271), (27553,-1.511039), (27554,-1.258761), (27555,-1.029709), (27556,-1.095610), (27557,-1.225612), (27558,-1.087600), (27559,-1.149786), (27560,-1.428426), (27561,-1.485037), (27562,-1.262023), (27563,-0.962832), (27564,-1.111878), (27565,-1.156877), (27566,-1.337973), (27567,-1.338381), (27568,-1.493930), (27569,-1.529639), (27570,-1.285258), (27571,-1.001395), (27572,-1.123500), (27573,-1.190330), (27574,-1.283637), (27575,-1.138194), (27576,-1.337405), (27577,-1.509211), (27578,-1.222097), (27579,-0.985148), (27580,-1.003206), (27581,-1.153646), (27582,-1.148015), (27583,-1.339794), (27584,-1.356924), (27585,-1.537091), (27586,-1.234648), (27587,-1.016279), (27588,-1.049201), (27589,-1.225188), (27590,-1.086712), (27591,-1.137749), (27592,-1.382946), (27593,-1.410759), (27594,-1.197964), (27595,-0.920139), (27596,-1.093338), (27597,-1.137873), (27598,-1.331975), (27599,-1.330990), (27600,-1.490254), (27601,-1.537576), (27602,-1.279260), (27603,-1.005152), (27604,-1.108212), (27605,-1.147173), (27606,-1.240480), (27607,-1.106184), (27608,-1.259875), (27609,-1.417747), (27610,-1.162217), (27611,-0.908083), (27612,-0.963765), (27613,-1.102127), (27614,-1.076988), (27615,-1.259942), (27616,-1.333276), (27617,-1.472567), (27618,-1.191955), (27619,-0.942465), (27620,-1.003722), (27621,-1.192714), (27622,-1.012433), (27623,-1.054646), (27624,-1.100109), (27625,-1.196667), (27626,-1.348965), (27627,-0.702331), (27628,-0.855558), (27629,-0.867578), (27630,-1.005012), (27631,-1.021212), (27632,-1.203702), (27633,-1.272855), (27634,-1.431655), (27635,-0.737643), (27636,-0.870432), (27637,-0.949339), (27638,-1.102565), (27639,-0.859114), (27640,-1.036958), (27641,-1.224557), (27642,-0.923508), (27643,-0.703281), (27644,-0.748280), (27645,-0.902436), (27646,-0.902843), (27647,-1.053747), (27648,-1.102927), (27649,-1.261262), (27650,-0.979257), (27651,-0.730232), (27652,-0.767799), (27653,-0.942856), (27654,-0.792768), (27655,-0.845664), (27656,-1.076461), (27657,-1.141898), (27658,-1.292801), (27659,-0.616905), (27660,-0.739010), (27661,-0.789119), (27662,-0.967428), (27663,-0.990596), (27664,-1.147539), (27665,-1.228304), (27666,-1.364344), (27667,-0.685661), (27668,-0.836564), (27669,-0.887137), (27670,-1.050118), (27671,-0.815956), (27672,-1.164270), (27673,-1.321213), (27674,-1.037814), (27675,-0.799007), (27676,-0.874663), (27677,-0.999555), (27678,-0.985099), (27679,-1.195923), (27680,-1.229309), (27681,-1.366279), (27682,-1.107963), (27683,-0.862653), (27684,-0.915549), (27685,-1.057627), (27686,-0.914970), (27687,-0.989233), (27688,-1.068140), (27689,-1.204180), (27690,-0.922175), (27691,-0.699626), (27692,-0.810119), (27693,-0.941049), (27694,-0.928451), (27695,-1.111405), (27696,-1.140147), (27697,-1.271542), (27698,-1.018336), (27699,-0.767452), (27700,-0.803161), (27701,-0.991689), (27702,-0.824879), (27703,-0.905644), (27704,-1.055154), (27705,-1.229284), (27706,-0.966787), (27707,-0.733090), (27708,-0.769264), (27709,-0.928064), (27710,-0.918717), (27711,-1.090058), (27712,-1.162928), (27713,-1.311045), (27714,-1.079205), (27715,-0.852939), (27716,-0.909551), (27717,-1.007502), (27718,-0.886677), (27719,-0.940501), (27720,-1.088618), (27721,-1.206079), (27722,-0.934758), (27723,-0.723356), (27724,-0.788792), (27725,-0.944806), (27726,-0.910841), (27727,-1.106336), (27728,-1.181063), (27729,-1.337541), (27730,-1.082941), (27731,-0.787930), (27732,-0.837110), (27733,-0.980582), (27734,-0.820739), (27735,-0.879209), (27736,-1.158313), (27737,-1.351950), (27738,-1.023960), (27739,-0.801411), (27740,-0.851055), (27741,-0.999636), (27742,-1.029772), (27743,-1.178353), (27744,-1.220101), (27745,-1.410952), (27746,-1.125695), (27747,-0.892926), (27748,-0.924920), (27749,-1.071179), (27750,-0.920625), (27751,-0.993959), (27752,-1.263774), (27753,-1.409104), (27754,-0.718344), (27755,-0.885040), (27756,-0.954658), (27757,-1.112994), (27758,-1.127336), (27759,-1.265699), (27760,-1.337174), (27761,-1.449989), (27762,-0.798711), (27763,-0.932893), (27764,-0.957919), (27765,-1.146912), (27766,-0.935974), (27767,-1.055757), (27768,-1.162999), (27769,-1.327373), (27770,-1.042581), (27771,-0.788445), (27772,-0.830657), (27773,-0.994103), (27774,-0.981505), (27775,-1.146344), (27776,-1.413372), (27777,-1.587500), (27778,-1.264620), (27779,-1.038818), (27780,-1.077779), (27781,-1.252836), (27782,-1.077665), (27783,-1.156572), (27784,-1.497920), (27785,-1.682731), (27786,-1.017054), (27787,-1.148913), (27788,-1.212028), (27789,-1.385227), (27790,-1.366126), (27791,-1.516566), (27792,-1.602441), (27793,-1.760312), (27794,-1.092777), (27795,-1.224172), (27796,-1.277532), (27797,-1.399637), (27798,-1.162688), (27799,-1.309411), (27800,-1.334438), (27801,-1.502064), (27802,-1.227026), (27803,-0.976142), (27804,-1.047617), (27805,-1.185051), (27806,-1.161305), (27807,-1.362838), (27808,-1.419450), (27809,-1.568496), (27810,-1.282775), (27811,-1.072303), (27812,-1.141456), (27813,-1.277496), (27814,-1.123226), (27815,-1.194702), (27816,-1.519791), (27817,-1.655367), (27818,-0.946027), (27819,-1.094144), (27820,-1.147968), (27821,-1.306769), (27822,-1.331794), (27823,-1.498027), (27824,-1.562535), (27825,-1.728767), (27826,-1.002706), (27827,-1.150823), (27828,-1.213472), (27829,-1.395033), (27830,-1.151116), (27831,-1.318277), (27832,-1.407868), (27833,-1.577352), (27834,-1.315320), (27835,-1.071404), (27836,-1.112687), (27837,-1.261269), (27838,-1.238916), (27839,-1.420941), (27840,-1.459438), (27841,-1.604767), (27842,-1.321833), (27843,-1.050048), (27844,-1.095511), (27845,-1.294722), (27846,-1.185974), (27847,-1.221683), (27848,-1.478492), (27849,-1.619641), (27850,-0.944674), (27851,-1.085359), (27852,-1.170305), (27853,-1.301235), (27854,-1.277954), (27855,-1.457656), (27856,-1.535635), (27857,-1.668888), (27858,-0.984166), (27859,-1.111381), (27860,-1.170315), (27861,-1.351875), (27862,-1.103779), (27863,-1.276978), (27864,-1.401406), (27865,-1.543020), (27866,-1.274485), (27867,-1.030104), (27868,-1.076033), (27869,-1.219505), (27870,-1.215732), (27871,-1.398221), (27872,-1.418138), (27873,-1.569506), (27874,-1.310726), (27875,-1.049624), (27876,-1.099268), (27877,-1.246455), (27878,-1.108444), (27879,-1.180848), (27880,-1.265329), (27881,-1.327050), (27882,-1.450549), (27883,-0.773724), (27884,-0.929272), (27885,-0.992387), (27886,-1.164193), (27887,-1.154382), (27888,-1.301570), (27889,-1.352143), (27890,-1.481680), (27891,-0.812287), (27892,-0.970159), (27893,-1.018873), (27894,-1.189751), (27895,-0.945834), (27896,-1.219365), (27897,-1.380488), (27898,-1.119385), (27899,-0.902409), (27900,-0.926506), (27901,-1.089487), (27902,-1.092217), (27903,-1.265416), (27904,-1.294623), (27905,-1.454817), (27906,-1.180708), (27907,-0.942366), (27908,-0.965533), (27909,-1.126657), (27910,-0.977497), (27911,-1.044792), (27912,-1.259331), (27913,-1.344277), (27914,-1.464989), (27915,-0.810460), (27916,-0.985517), (27917,-1.047238), (27918,-1.192568), (27919,-1.208769), (27920,-1.359673), (27921,-1.388879), (27922,-1.524455), (27923,-0.896866), (27924,-1.048698), (27925,-1.093233), (27926,-1.273865), (27927,-1.038309), (27928,-1.431679), (27929,-1.182653), (27930,-1.323803), (27931,-0.947041), (27932,-1.084010), (27933,-1.068625), (27934,-1.219064), (27935,-1.346279), (27936,-1.453520), (27937,-1.167800), (27938,-1.317775), (27939,-1.003719), (27940,-1.152301), (27941,-1.002677), (27942,-1.127104), (27943,-1.076882), (27944,-1.174369), (27945,-1.343854), (27946,-1.039088), (27947,-0.797959), (27948,-0.808121), (27949,-0.978533), (27950,-0.935279), (27951,-1.142386), (27952,-1.193889), (27953,-1.362908), (27954,-1.082296), (27955,-0.866249), (27956,-0.864799), (27957,-1.049611), (27958,-0.890233), (27959,-0.983075), (27960,-1.348111), (27961,-1.034056), (27962,-1.181708), (27963,-0.808662), (27964,-0.952134), (27965,-0.971586), (27966,-1.130851), (27967,-1.237628), (27968,-1.384352), (27969,-1.088876), (27970,-1.233277), (27971,-0.912255), (27972,-1.049224), (27973,-0.915857), (27974,-1.071406), (27975,-1.036048), (27976,-1.199957), (27977,-1.404743), (27978,-1.135743), (27979,-0.883930), (27980,-0.927072), (27981,-1.081691), (27982,-1.039830), (27983,-1.233003), (27984,-1.288221), (27985,-1.447486), (27986,-1.166410), (27987,-0.928997), (27988,-0.974461), (27989,-1.146267), (27990,-0.968773), (27991,-1.056505), (27992,-1.306812), (27993,-0.994614), (27994,-1.153415), (27995,-0.833321), (27996,-0.978187), (27997,-0.967911), (27998,-1.134143), (27999,-1.202832), (28000,-1.367671), (28001,-1.089846), (28002,-1.257007), (28003,-0.929017), (28004,-1.031614), (28005,-0.868055), (28006,-1.040790), (28007,-0.985458), (28008,-1.263634), (28009,-1.409892), (28010,-0.740499), (28011,-0.909518), (28012,-0.994000), (28013,-1.142117), (28014,-1.157388), (28015,-1.298537), (28016,-1.348182), (28017,-1.481435), (28018,-0.846879), (28019,-0.986634), (28020,-1.032098), (28021,-1.176964), (28022,-0.939086), (28023,-1.121576), (28024,-1.180509), (28025,-1.330949), (28026,-1.068453), (28027,-0.825000), (28028,-0.882541), (28029,-1.039948), (28030,-1.037569), (28031,-1.220523), (28032,-1.512169), (28033,-1.650067), (28034,-1.352733), (28035,-1.144583), (28036,-1.217452), (28037,-1.359995), (28038,-1.220126), (28039,-1.273950), (28040,-1.347748), (28041,-1.497722), (28042,-1.215718), (28043,-0.975982), (28044,-1.053496), (28045,-1.191858), (28046,-1.182047), (28047,-1.340383), (28048,-1.408607), (28049,-1.563226), (28050,-1.275183), (28051,-1.034518), (28052,-1.090201), (28053,-1.253182), (28054,-1.117028), (28055,-1.151808), (28056,-1.437880), (28057,-1.597145), (28058,-1.291915), (28059,-1.054037), (28060,-1.104145), (28061,-1.274094), (28062,-1.283327), (28063,-1.448165), (28064,-1.497810), (28065,-1.666829), (28066,-1.329549), (28067,-1.113503), (28068,-1.168721), (28069,-1.333095), (28070,-1.154208), (28071,-1.219180), (28072,-1.262786), (28073,-1.341228), (28074,-1.513964), (28075,-0.845499), (28076,-0.990830), (28077,-1.058124), (28078,-1.204848), (28079,-1.217797), (28080,-1.365914), (28081,-1.430422), (28082,-1.618485), (28083,-0.940266), (28084,-1.092099), (28085,-1.148246), (28086,-1.271745), (28087,-1.076136), (28088,-1.460217), (28089,-1.638061), (28090,-1.361630), (28091,-1.116784), (28092,-1.142275), (28093,-1.306185), (28094,-1.293122), (28095,-1.518345), (28096,-1.557770), (28097,-1.697991), (28098,-1.418773), (28099,-1.181359), (28100,-1.216604), (28101,-1.364721), (28102,-1.196982), (28103,-1.235942), (28104,-1.248892), (28105,-1.318045), (28106,-1.463839), (28107,-0.800949), (28108,-0.981580), (28109,-1.027508), (28110,-1.179805), (28111,-1.163027), (28112,-1.333904), (28113,-1.396554), (28114,-1.569289), (28115,-0.870168), (28116,-1.042439), (28117,-1.103696), (28118,-1.257851), (28119,-1.035766), (28120,-1.423097), (28121,-1.623238), (28122,-1.329620), (28123,-1.082452), (28124,-1.129309), (28125,-1.290432), (28126,-1.256003), (28127,-1.428274), (28128,-1.511361), (28129,-1.649724), (28130,-1.382583), (28131,-1.136809), (28132,-1.166014), (28133,-1.335963), (28134,-1.177978), (28135,-1.255957), (28136,-1.325573), (28137,-1.361283), (28138,-1.540985), (28139,-0.848832), (28140,-0.995555), (28141,-1.046593), (28142,-1.189601), (28143,-1.210446), (28144,-1.354847), (28145,-1.437006), (28146,-1.565614), (28147,-0.872996), (28148,-1.035977), (28149,-1.113490), (28150,-1.300160), (28151,-1.099442), (28152,-1.156983), (28153,-1.284197), (28154,-0.980825), (28155,-1.170747), (28156,-0.799094), (28157,-0.946282), (28158,-0.944832), (28159,-1.073905), (28160,-1.180682), (28161,-1.332980), (28162,-1.034252), (28163,-1.183763), (28164,-0.859953), (28165,-1.002496), (28166,-0.860304), (28167,-1.044187), (28168,-1.151429), (28169,-1.208040), (28170,-1.378918), (28171,-1.077404), (28172,-0.839990), (28173,-0.881273), (28174,-1.039609), (28175,-1.047449), (28176,-1.193708), (28177,-1.259609), (28178,-1.436525), (28179,-1.136404), (28180,-0.930113), (28181,-0.971860), (28182,-1.111616), (28183,-0.974534), (28184,-1.132870), (28185,-1.320468), (28186,-1.045895), (28187,-1.201444), (28188,-0.846049), (28189,-0.995095), (28190,-0.984355), (28191,-1.138510), (28192,-1.241571), (28193,-1.394797), (28194,-1.112328), (28195,-1.227930), (28196,-0.889721), (28197,-1.055025), (28198,-0.932341), (28199,-1.102290), (28200,-1.300572), (28201,-1.440328), (28202,-1.138815), (28203,-0.901401), (28204,-0.947793), (28205,-1.116348), (28206,-1.113969), (28207,-1.276950), (28208,-1.315446), (28209,-1.514193), (28210,-1.255412), (28211,-1.015212), (28212,-1.056960), (28213,-1.184175), (28214,-1.066136), (28215,-1.136218), (28216,-1.149632), (28217,-1.306574), (28218,-1.038504), (28219,-1.192659), (28220,-0.834941), (28221,-1.015573), (28222,-0.997401), (28223,-1.147840), (28224,-1.227212), (28225,-1.378581), (28226,-1.131878), (28227,-1.256770), (28228,-0.910664), (28229,-1.106160), (28230,-0.956536), (28231,-1.121839), (28232,-1.149652), (28233,-1.300556), (28234,-1.018086), (28235,-1.162023), (28236,-0.814524), (28237,-0.978434), (28238,-1.034581), (28239,-1.182698), (28240,-1.260676), (28241,-1.400433), (28242,-1.157910), (28243,-1.279086), (28244,-0.932981), (28245,-1.082491), (28246,-0.917074), (28247,-1.084700), (28248,-1.189619), (28249,-1.332162), (28250,-1.035293), (28251,-1.194558), (28252,-0.851239), (28253,-1.015614), (28254,-1.004874), (28255,-1.142772), (28256,-1.210531), (28257,-1.368403), (28258,-1.105906), (28259,-1.196890), (28260,-0.880513), (28261,-1.026772), (28262,-0.887831), (28263,-1.030838), (28264,-1.203574), (28265,-1.345653), (28266,-1.094769), (28267,-0.852710), (28268,-0.897709), (28269,-1.056509), (28270,-1.035086), (28271,-1.187383), (28272,-1.292303), (28273,-1.484082), (28274,-1.198825), (28275,-0.968844), (28276,-1.031494), (28277,-1.173108), (28278,-0.957061), (28279,-1.003919), (28280,-1.344336), (28281,-1.502672), (28282,-1.221132), (28283,-0.954455), (28284,-1.005028), (28285,-1.174047), (28286,-1.154946), (28287,-1.320249), (28288,-1.410304), (28289,-1.554706), (28290,-1.284777), (28291,-1.048757), (28292,-1.106298), (28293,-1.258131), (28294,-1.093643), (28295,-1.162796), (28296,-1.513897), (28297,-1.540781), (28298,-1.288968), (28299,-1.009750), (28300,-1.158332), (28301,-1.198686), (28302,-1.370492), (28303,-1.356964), (28304,-1.510656), (28305,-1.585383), (28306,-1.338215), (28307,-1.023231), (28308,-1.190856), (28309,-1.254900), (28310,-1.333343), (28311,-1.196260), (28312,-1.330907), (28313,-1.386124), (28314,-1.543995), (28315,-0.878782), (28316,-1.015752), (28317,-1.074221), (28318,-1.242311), (28319,-1.234358), (28320,-1.384797), (28321,-1.469279), (28322,-1.615073), (28323,-0.910843), (28324,-1.085901), (28325,-1.107675), (28326,-1.260437), (28327,-1.026275), (28328,-1.484210), (28329,-1.508771), (28330,-1.254171), (28331,-1.003287), (28332,-1.128180), (28333,-1.195475), (28334,-1.396544), (28335,-1.384411), (28336,-1.585479), (28337,-1.622583), (28338,-1.351261), (28339,-1.064146), (28340,-1.227592), (28341,-1.282810), (28342,-1.353356), (28343,-1.213486), (28344,-1.356958), (28345,-1.452587), (28346,-1.567725), (28347,-0.899261), (28348,-1.038552), (28349,-1.102596), (28350,-1.254429), (28351,-1.246940), (28352,-1.384838), (28353,-1.462816), (28354,-1.635087), (28355,-0.966623), (28356,-1.104986), (28357,-1.196898), (28358,-1.332938), (28359,-1.093203), (28360,-1.412718), (28361,-1.443783), (28362,-1.236097), (28363,-0.955485), (28364,-1.108712), (28365,-1.136989), (28366,-1.316227), (28367,-1.315706), (28368,-1.497731), (28369,-1.529724), (28370,-1.311819), (28371,-1.045608), (28372,-1.225774), (28373,-1.280063), (28374,-1.351538), (28375,-1.226069), (28376,-1.342600), (28377,-1.408966), (28378,-1.584953), (28379,-0.893263), (28380,-1.015833), (28381,-1.057116), (28382,-1.214988), (28383,-1.212144), (28384,-1.403459), (28385,-1.434058), (28386,-1.598433), (28387,-0.912782), (28388,-1.079943), (28389,-1.155599), (28390,-1.296284), (28391,-1.059800), (28392,-1.206988), (28393,-1.249665), (28394,-1.432154), (28395,-0.775302), (28396,-0.922954), (28397,-0.993500), (28398,-1.127683), (28399,-1.179650), (28400,-1.293858), (28401,-1.372301), (28402,-1.498122), (28403,-0.808755), (28404,-0.976381), (28405,-1.040889), (28406,-1.171820), (28407,-0.939980), (28408,-1.219085), (28409,-1.291954), (28410,-1.427065), (28411,-0.732124), (28412,-0.902073), (28413,-0.971225), (28414,-1.110053), (28415,-1.112782), (28416,-1.246965), (28417,-1.301253), (28418,-1.466092), (28419,-0.753501), (28420,-0.948532), (28421,-1.001427), (28422,-1.158370), (28423,-0.923279), (28424,-1.224214), (28425,-1.280826), (28426,-1.442878), (28427,-0.738183), (28428,-0.911383), (28429,-0.979606), (28430,-1.123078), (28431,-1.162503), (28432,-1.330129), (28433,-1.356084), (28434,-1.508382), (28435,-0.844562), (28436,-0.985712), (28437,-1.051149), (28438,-1.176505), (28439,-0.914473), (28440,-1.207978), (28441,-1.393719), (28442,-1.125648), (28443,-0.878016), (28444,-0.908151), (28445,-1.075313), (28446,-1.070146), (28447,-1.229876), (28448,-1.296706), (28449,-1.480589), (28450,-1.206016), (28451,-0.948629), (28452,-0.964366), (28453,-1.120843), (28454,-0.989334), (28455,-1.037121), (28456,-1.125782), (28457,-1.283189), (28458,-0.996539), (28459,-0.757732), (28460,-0.793442), (28461,-0.965248), (28462,-0.953114), (28463,-1.136533), (28464,-1.160165), (28465,-1.340332), (28466,-1.062972), (28467,-0.844603), (28468,-0.897498), (28469,-1.052583), (28470,-0.892276), (28471,-0.947493), (28472,-1.214986), (28473,-1.419771), (28474,-1.128012), (28475,-0.900352), (28476,-0.945816), (28477,-1.122732), (28478,-1.107346), (28479,-1.276830), (28480,-1.357595), (28481,-1.528008), (28482,-1.246932), (28483,-0.983507), (28484,-1.012713), (28485,-1.225395), (28486,-1.056262), (28487,-1.125880), (28488,-1.230334), (28489,-1.385883), (28490,-1.112703), (28491,-0.885509), (28492,-0.890097), (28493,-1.037285), (28494,-1.006571), (28495,-1.200209), (28496,-1.240563), (28497,-1.407260), (28498,-1.124326), (28499,-0.900847), (28500,-0.971858), (28501,-1.117188), (28502,-0.950378), (28503,-1.023246), (28504,-1.201091), (28505,-1.355711), (28506,-1.064416), (28507,-0.830254), (28508,-0.888724), (28509,-1.071213), (28510,-1.051648), (28511,-1.231815), (28512,-1.275420), (28513,-1.433292), (28514,-1.150358), (28515,-0.910622), (28516,-0.944009), (28517,-1.091661), (28518,-0.944824), (28519,-1.025125), (28520,-1.269392), (28521,-1.317643), (28522,-1.083481), (28523,-0.791722), (28524,-0.945412), (28525,-0.988089), (28526,-1.154786), (28527,-1.162161), (28528,-1.333503), (28529,-1.371070), (28530,-1.154559), (28531,-0.853509), (28532,-1.043431), (28533,-1.109797), (28534,-1.141790), (28535,-1.011210), (28536,-1.176514), (28537,-1.306980), (28538,-1.055631), (28539,-0.797780), (28540,-0.874365), (28541,-0.982071), (28542,-0.970402), (28543,-1.163110), (28544,-1.074799), (28545,-1.126766), (28546,-0.908861), (28547,-0.625927), (28548,-0.761039), (28549,-0.809753), (28550,-0.867294), (28551,-0.705129), (28552,-0.957292), (28553,-0.978602), (28554,-0.756982), (28555,-0.476835), (28556,-0.654680), (28557,-0.725690), (28558,-0.902606), (28559,-0.881182), (28560,-1.039518), (28561,-1.102168), (28562,-0.855001), (28563,-0.559990), (28564,-0.723899), (28565,-0.774937), (28566,-0.905403), (28567,-0.697717), (28568,-0.960100), (28569,-1.021356), (28570,-0.793697), (28571,-0.546994), (28572,-0.709046), (28573,-0.772160), (28574,-0.949540), (28575,-0.914182), (28576,-1.083665), (28577,-1.114730), (28578,-0.833189), (28579,-0.535856), (28580,-0.682579), (28581,-0.754519), (28582,-0.836678), (28583,-0.697738), (28584,-1.093430), (28585,-0.797955), (28586,-0.960471), (28587,-0.694259), (28588,-0.824260), (28589,-0.869260), (28590,-0.979752), (28591,-1.025681), (28592,-1.187268), (28593,-0.840698), (28594,-0.947939), (28595,-0.742112), (28596,-0.847495), (28597,-0.830717), (28598,-0.975582), (28599,-0.817597), (28600,-1.026563), (28601,-1.062737), (28602,-0.834148), (28603,-0.564220), (28604,-0.714660), (28605,-0.781955), (28606,-0.994637), (28607,-0.985290), (28608,-1.137587), (28609,-1.140782), (28610,-0.899188), (28611,-0.629724), (28612,-0.774126), (28613,-0.826092), (28614,-0.893852), (28615,-0.736795), (28616,-0.890951), (28617,-0.954065), (28618,-0.767746), (28619,-0.501534), (28620,-0.669160), (28621,-0.722984), (28622,-0.873423), (28623,-0.848749), (28624,-1.020555), (28625,-1.079024), (28626,-0.887596), (28627,-0.598159), (28628,-0.735593), (28629,-0.781521), (28630,-0.825126), (28631,-0.652278), (28632,-0.999663), (28633,-1.066029), (28634,-0.821183), (28635,-0.554507), (28636,-0.689153), (28637,-0.750875), (28638,-0.951015), (28639,-0.948171), (28640,-1.069347), (28641,-1.103198), (28642,-0.857889), (28643,-0.599573), (28644,-0.764411), (28645,-0.830778), (28646,-0.878099), (28647,-0.724759), (28648,-0.790660), (28649,-0.927165), (28650,-0.604749), (28651,-0.734751), (28652,-0.465287), (28653,-0.627804), (28654,-0.711820), (28655,-0.843680), (28656,-0.819470), (28657,-0.999636), (28658,-0.671646), (28659,-0.798397), (28660,-0.513605), (28661,-0.666367), (28662,-0.641227), (28663,-0.761010), (28664,-0.895657), (28665,-0.930901), (28666,-0.710210), (28667,-0.421237), (28668,-0.619520), (28669,-0.686815), (28670,-0.851189), (28671,-0.820011), (28672,-0.940258), (28673,-1.004302), (28674,-0.768282), (28675,-0.484883), (28676,-0.653438), (28677,-0.734668), (28678,-0.791744), (28679,-0.589167), (28680,-0.773050), (28681,-0.962507), (28682,-0.613615), (28683,-0.790996), (28684,-0.520602), (28685,-0.659429), (28686,-0.744376), (28687,-0.892957), (28688,-0.890113), (28689,-1.034514), (28690,-0.701879), (28691,-0.843958), (28692,-0.565669), (28693,-0.730043), (28694,-0.684930), (28695,-0.840944), (28696,-0.787005), (28697,-0.937445), (28698,-0.651260), (28699,-0.393408), (28700,-0.443981), (28701,-0.615323), (28702,-0.592971), (28703,-0.771279), (28704,-0.814421), (28705,-1.005271), (28706,-0.666598), (28707,-0.422682), (28708,-0.496015), (28709,-0.618585), (28710,-0.464780), (28711,-0.533933), (28712,-0.792600), (28713,-0.838528), (28714,-0.634558), (28715,-0.359056), (28716,-0.511818), (28717,-0.559139), (28718,-0.735590), (28719,-0.697910), (28720,-0.852065), (28721,-0.933759), (28722,-0.694023), (28723,-0.424560), (28724,-0.589399), (28725,-0.637185), (28726,-0.678932), (28727,-0.546495), (28728,-0.908744), (28729,-1.061505), (28730,-0.344734), (28731,-0.485419), (28732,-0.546675), (28733,-0.685502), (28734,-0.722605), (28735,-0.888373), (28736,-0.913399), (28737,-1.088921), (28738,-0.416740), (28739,-0.593191), (28740,-0.643765), (28741,-0.792811), (28742,-0.573512), (28743,-0.716520), (28744,-0.890649), (28745,-0.889198), (28746,-0.686158), (28747,-0.397649), (28748,-0.570385), (28749,-0.618171), (28750,-0.815989), (28751,-0.784346), (28752,-0.934786), (28753,-0.989075), (28754,-0.761416), (28755,-0.458973), (28756,-0.619167), (28757,-0.673456), (28758,-0.715668), (28759,-0.548858), (28760,-0.641700), (28761,-0.795391), (28762,-0.522211), (28763,-0.319635), (28764,-0.368350), (28765,-0.542014), (28766,-0.546138), (28767,-0.699829), (28768,-0.748079), (28769,-0.942181), (28770,-0.651815), (28771,-0.438556), (28772,-0.465439), (28773,-0.613092), (28774,-0.481119), (28775,-0.566994), (28776,-0.917630), (28777,-0.608220), (28778,-0.776775), (28779,-0.472009), (28780,-0.601547), (28781,-0.690208), (28782,-0.838325), (28783,-0.805289), (28784,-1.010539), (28785,-0.655144), (28786,-0.796758), (28787,-0.534726), (28788,-0.694920), (28789,-0.676283), (28790,-0.796531), (28791,-0.652481), (28792,-0.868414), (28793,-0.889259), (28794,-0.658813), (28795,-0.384704), (28796,-0.556046), (28797,-0.609406), (28798,-0.786786), (28799,-0.747248), (28800,-0.937634), (28801,-1.084357), (28802,-0.554312), (28803,-0.691745), (28804,-0.776227), (28805,-0.895545), (28806,-0.554085), (28807,-0.709634), (28808,-0.868899), (28809,-1.031879), (28810,-0.621674), (28811,-0.725199), (28812,-0.795746), (28813,-0.959656), (28814,-0.699482), (28815,-0.837380), (28816,-0.898172), (28817,-1.057437), (28818,-0.506489), (28819,-0.653213), (28820,-0.682419), (28821,-0.809634), (28822,-0.447736), (28823,-0.622794), (28824,-0.848945), (28825,-0.933891), (28826,-0.702981), (28827,-0.650901), (28828,-0.819920), (28829,-0.899292), (28830,-1.049266), (28831,-0.767726), (28832,-0.950215), (28833,-0.980351), (28834,-0.748511), (28835,-0.613751), (28836,-0.730282), (28837,-0.765062), (28838,-0.841183), (28839,-0.596338), (28840,-0.818309), (28841,-0.870276), (28842,-0.612889), (28843,-0.589143), (28844,-0.737724), (28845,-0.828709), (28846,-0.997728), (28847,-0.726406), (28848,-0.893568), (28849,-0.934851), (28850,-0.712765), (28851,-0.577541), (28852,-0.751205), (28853,-0.798991), (28854,-0.838416), (28855,-0.565237), (28856,-0.875927), (28857,-0.933932), (28858,-0.700699), (28859,-0.723402), (28860,-0.866410), (28861,-0.916983), (28862,-1.088789), (28863,-0.810036), (28864,-0.984164), (28865,-1.059355), (28866,-0.793608), (28867,-0.633300), (28868,-0.808823), (28869,-0.846854), (28870,-0.909505), (28871,-0.627964), (28872,-0.834143), (28873,-0.860562), (28874,-0.632903), (28875,-0.610550), (28876,-0.797220), (28877,-0.843613), (28878,-1.024245), (28879,-0.700900), (28880,-0.864810), (28881,-0.926531), (28882,-0.689582), (28883,-0.520913), (28884,-0.666243), (28885,-0.741899), (28886,-0.816625), (28887,-0.542982), (28888,-0.915914), (28889,-0.991105), (28890,-0.814541), (28891,-0.798227), (28892,-0.929157), (28893,-0.983446), (28894,-1.162684), (28895,-0.887182), (28896,-1.045983), (28897,-1.096555), (28898,-0.835917), (28899,-0.684900), (28900,-0.832553), (28901,-0.838069), (28902,-0.940201), (28903,-0.630327), (28904,-0.818390), (28905,-0.869893), (28906,-0.655239), (28907,-0.630100), (28908,-0.775894), (28909,-0.813461), (28910,-1.003383), (28911,-0.728810), (28912,-0.869959), (28913,-0.925177), (28914,-0.678474), (28915,-0.536746), (28916,-0.671858), (28917,-0.745191), (28918,-0.830601), (28919,-0.573679), (28920,-0.619142), (28921,-0.650207), (28922,-0.805291), (28923,-0.415523), (28924,-0.564105), (28925,-0.602601), (28926,-0.767440), (28927,-0.521666), (28928,-0.747353), (28929,-0.799784), (28930,-0.954404), (28931,-0.376051), (28932,-0.531136), (28933,-0.598895), (28934,-0.737258), (28935,-0.359567), (28936,-0.669793), (28937,-0.720830), (28938,-0.885669), (28939,-0.493115), (28940,-0.694184), (28941,-0.721532), (28942,-0.875223), (28943,-0.636416), (28944,-0.755735), (28945,-0.811881), (28946,-0.931200), (28947,-0.401155), (28948,-0.552987), (28949,-0.599380), (28950,-0.751678), (28951,-0.380025), (28952,-0.636369), (28953,-0.805388), (28954,-0.813693), (28955,-0.581853), (28956,-0.664941), (28957,-0.791691), (28958,-0.500861), (28959,-0.644333), (28960,-0.678649), (28961,-0.853706), (28962,-0.716624), (28963,-0.473171), (28964,-0.546969), (28965,-0.693228), (28966,-0.405649), (28967,-0.462261), (28968,-0.848664), (28969,-1.007464), (28970,-0.621412), (28971,-0.730047), (28972,-0.818244), (28973,-0.974258), (28974,-0.739631), (28975,-0.888213), (28976,-0.945753), (28977,-1.068323), (28978,-0.577296), (28979,-0.727735), (28980,-0.789456), (28981,-0.933393), (28982,-0.560346), (28983,-0.699638), (28984,-0.690291), (28985,-0.835621), (28986,-0.816985), (28987,-0.605583), (28988,-0.645937), (28989,-0.810312), (28990,-0.501366), (28991,-0.671778), (28992,-0.746505), (28993,-0.913202), (28994,-0.767758), (28995,-0.550783), (28996,-0.609717), (28997,-0.752260), (28998,-0.438204), (28999,-0.507357), (29000,-0.694027), (29001,-0.840751), (29002,-0.840694), (29003,-0.589811), (29004,-0.631093), (29005,-0.781533), (29006,-0.494883), (29007,-0.651825), (29008,-0.721443), (29009,-0.872811), (29010,-0.706465), (29011,-0.486238), (29012,-0.532631), (29013,-0.687251), (29014,-0.435438), (29015,-0.492978), (29016,-0.624838), (29017,-0.800360), (29018,-0.800768), (29019,-0.560103), (29020,-0.597206), (29021,-0.784805), (29022,-0.477717), (29023,-0.635124), (29024,-0.686626), (29025,-0.865864), (29026,-0.736213), (29027,-0.522489), (29028,-0.550302), (29029,-0.707245), (29030,-0.428026), (29031,-0.486961), (29032,-0.750272), (29033,-0.883061), (29034,-0.522092), (29035,-0.662312), (29036,-0.717066), (29037,-0.867505), (29038,-0.607331), (29039,-0.759164), (29040,-0.820421), (29041,-0.936952), (29042,-0.410623), (29043,-0.559205), (29044,-0.639505), (29045,-0.786229), (29046,-0.428046), (29047,-0.571983), (29048,-0.844120), (29049,-0.964368), (29050,-0.547659), (29051,-0.702743), (29052,-0.731021), (29053,-0.890750), (29054,-0.649621), (29055,-0.774048), (29056,-0.999272), (29057,-1.087469), (29058,-0.835191), (29059,-0.688354), (29060,-0.844367), (29061,-0.899121), (29062,-0.976170), (29063,-0.710887), (29064,-0.890590), (29065,-0.981574), (29066,-0.729297), (29067,-0.725060), (29068,-0.853203), (29069,-0.930253), (29070,-1.078834), (29071,-0.810763), (29072,-0.961203), (29073,-1.003416), (29074,-0.762750), (29075,-0.613127), (29076,-0.749167), (29077,-0.828074), (29078,-0.897691), (29079,-0.583172), (29080,-0.933808), (29081,-0.972304), (29082,-0.706557), (29083,-0.706964), (29084,-0.861584), (29085,-0.897758), (29086,-1.113691), (29087,-0.823325), (29088,-1.001634), (29089,-1.036880), (29090,-0.800395), (29091,-0.611753), (29092,-0.803068), (29093,-0.872221), (29094,-0.924187), (29095,-0.662156), (29096,-0.735025), (29097,-0.882213), (29098,-0.545862), (29099,-0.721849), (29100,-0.727366), (29101,-0.894991), (29102,-0.955784), (29103,-1.110868), (29104,-0.838153), (29105,-0.985805), (29106,-0.649919), (29107,-0.799894), (29108,-0.607072), (29109,-0.779807), (29110,-0.747700), (29111,-0.903714), (29112,-0.886470), (29113,-1.047129), (29114,-0.678263), (29115,-0.839850), (29116,-0.834219), (29117,-0.991627), (29118,-1.057528), (29119,-1.240946), (29120,-0.967302), (29121,-1.120529), (29122,-0.754915), (29123,-0.902103), (29124,-0.791032), (29125,-0.944258), (29126,-0.919119), (29127,-1.042618), (29128,-0.706731), (29129,-0.882253), (29130,-0.541722), (29131,-0.676368), (29132,-0.671202), (29133,-0.816068), (29134,-0.905658), (29135,-1.067710), (29136,-0.769913), (29137,-0.946828), (29138,-0.583537), (29139,-0.743731), (29140,-0.584817), (29141,-0.731540), (29142,-0.685034), (29143,-0.822932), (29144,-0.840061), (29145,-1.001184), (29146,-0.648576), (29147,-0.799480), (29148,-0.811964), (29149,-0.945218), (29150,-1.032021), (29151,-1.175029), (29152,-0.912997), (29153,-1.064366), (29154,-0.750775), (29155,-0.881241), (29156,-0.751126), (29157,-0.886702), (29158,-0.862491), (29159,-1.020827), (29160,-0.758795), (29161,-0.931530), (29162,-0.578458), (29163,-0.718678), (29164,-0.720015), (29165,-0.872777), (29166,-0.938214), (29167,-1.094227), (29168,-0.814545), (29169,-1.004466), (29170,-0.642104), (29171,-0.808800), (29172,-0.646635), (29173,-0.777566), (29174,-0.717589), (29175,-0.890324), (29176,-0.463861), (29177,-0.612443), (29178,-0.666267), (29179,-0.440466), (29180,-0.446913), (29181,-0.620577), (29182,-0.651641), (29183,-0.824840), (29184,-0.610652), (29185,-0.730899), (29186,-0.806090), (29187,-0.560316), (29188,-0.377248), (29189,-0.519327), (29190,-0.588015), (29191,-0.650201), (29192,-0.516370), (29193,-0.658448), (29194,-0.723420), (29195,-0.481827), (29196,-0.455294), (29197,-0.617810), (29198,-0.657235), (29199,-0.875491), (29200,-0.592557), (29201,-0.753680), (29202,-0.807040), (29203,-0.550582), (29204,-0.434401), (29205,-0.594131), (29206,-0.627053), (29207,-0.692025), (29208,-0.629726), (29209,-0.699344), (29210,-0.849783), (29211,-0.446081), (29212,-0.573760), (29213,-0.655454), (29214,-0.816577), (29215,-0.571267), (29216,-0.715668), (29217,-0.801543), (29218,-0.937118), (29219,-0.409860), (29220,-0.564016), (29221,-0.611802), (29222,-0.739945), (29223,-0.373867), (29224,-0.800681), (29225,-0.821062), (29226,-0.600370), (29227,-0.604493), (29228,-0.745179), (29229,-0.823157), (29230,-0.980099), (29231,-0.690198), (29232,-0.842496), (29233,-0.873560), (29234,-0.636611), (29235,-0.488380), (29236,-0.662973), (29237,-0.704721), (29238,-0.759475), (29239,-0.510449), (29240,-0.630232), (29241,-0.684056), (29242,-0.824276), (29243,-0.428471), (29244,-0.569620), (29245,-0.640166), (29246,-0.803147), (29247,-0.569914), (29248,-0.700380), (29249,-0.751418), (29250,-0.893961), (29251,-0.382031), (29252,-0.512497), (29253,-0.559354), (29254,-0.720013), (29255,-0.361366), (29256,-0.598202), (29257,-0.666890), (29258,-0.818259), (29259,-0.411769), (29260,-0.602620), (29261,-0.648548), (29262,-0.783659), (29263,-0.518840), (29264,-0.676712), (29265,-0.741684), (29266,-0.906058), (29267,-0.366723), (29268,-0.540387), (29269,-0.573774), (29270,-0.724213), (29271,-0.359993), (29272,-0.614015), (29273,-0.680380), (29274,-0.879127), (29275,-0.434550), (29276,-0.617039), (29277,-0.653677), (29278,-0.797149), (29279,-0.540227), (29280,-0.712962), (29281,-0.757497), (29282,-0.926052), (29283,-0.376962), (29284,-0.509286), (29285,-0.576581), (29286,-0.726556), (29287,-0.390206), (29288,-0.733875), (29289,-0.771906), (29290,-0.533564), (29291,-0.487987), (29292,-0.667689), (29293,-0.726159), (29294,-0.932802), (29295,-0.636862), (29296,-0.822603), (29297,-0.850416), (29298,-0.599532), (29299,-0.450373), (29300,-0.613353), (29301,-0.668107), (29302,-0.753053), (29303,-0.426921), (29304,-0.840729), (29305,-0.917313), (29306,-0.680364), (29307,-0.655225), (29308,-0.830283), (29309,-0.847877), (29310,-1.049875), (29311,-0.758116), (29312,-1.104572), (29313,-1.152822), (29314,-0.902867), (29315,-0.753244), (29316,-0.893464), (29317,-0.943108), (29318,-1.036415), (29319,-0.756268), (29320,-1.012147), (29321,-1.053895), (29322,-0.769103), (29323,-0.788555), (29324,-0.955717), (29325,-1.042985), (29326,-1.220829), (29327,-0.923961), (29328,-1.086477), (29329,-1.120792), (29330,-0.918216), (29331,-0.773237), (29332,-0.897201), (29333,-0.970069), (29334,-1.047583), (29335,-0.787874), (29336,-0.757160), (29337,-0.911315), (29338,-0.921013), (29339,-0.701251), (29340,-0.688652), (29341,-0.867890), (29342,-0.902206), (29343,-1.128823), (29344,-0.837528), (29345,-0.986574), (29346,-1.040399), (29347,-0.769541), (29348,-0.632923), (29349,-0.796833), (29350,-0.840903), (29351,-0.908198), (29352,-0.829178), (29353,-0.983797), (29354,-0.641408), (29355,-0.792777), (29356,-0.787146), (29357,-0.955236), (29358,-1.018350), (29359,-1.179937), (29360,-0.884927), (29361,-1.047443), (29362,-0.689725), (29363,-0.849919), (29364,-0.690541), (29365,-0.852128), (29366,-0.821415), (29367,-0.991827), (29368,-0.944392), (29369,-1.085077), (29370,-0.741294), (29371,-0.903346), (29372,-0.891212), (29373,-1.024930), (29374,-1.114986), (29375,-1.265889), (29376,-0.990387), (29377,-1.160335), (29378,-0.787289), (29379,-0.955844), (29380,-0.846166), (29381,-0.977562), (29382,-0.947778), (29383,-1.109365), (29384,-0.885422), (29385,-1.049331), (29386,-0.694865), (29387,-0.844840), (29388,-0.845712), (29389,-0.965960), (29390,-1.046260), (29391,-1.184623), (29392,-0.931417), (29393,-1.069779), (29394,-0.729248), (29395,-0.869004), (29396,-0.736102), (29397,-0.892115), (29398,-0.861867), (29399,-1.038318), (29400,-0.771176), (29401,-0.965278), (29402,-0.984266), (29403,-0.729666), (29404,-0.731003), (29405,-0.913492), (29406,-0.961743), (29407,-1.144697), (29408,-0.842719), (29409,-1.029853), (29410,-1.076246), (29411,-0.827220), (29412,-0.681312), (29413,-0.841506), (29414,-0.869783), (29415,-0.907350), (29416,-0.625810), (29417,-0.791578), (29418,-0.857014), (29419,-0.625175), (29420,-0.639517), (29421,-0.817826), (29422,-0.830776), (29423,-1.013265), (29424,-0.739157), (29425,-0.916072), (29426,-0.980116), (29427,-0.697646), (29428,-0.518294), (29429,-0.696603), (29430,-0.762041), (29431,-0.820046), (29432,-0.567304), (29433,-0.735394), (29434,-0.795257), (29435,-0.550876), (29436,-0.512731), (29437,-0.695685), (29438,-0.747187), (29439,-0.936180), (29440,-0.604009), (29441,-0.736333), (29442,-0.793874), (29443,-0.544383), (29444,-0.405443), (29445,-0.556811), (29446,-0.632002), (29447,-0.731812), (29448,-0.643036), (29449,-0.786973), (29450,-0.839404), (29451,-0.574586), (29452,-0.585212), (29453,-0.751445), (29454,-0.782509), (29455,-0.958495), (29456,-0.665343), (29457,-0.816711), (29458,-0.858459), (29459,-0.635909), (29460,-0.506258), (29461,-0.659485), (29462,-0.721670), (29463,-0.790359), (29464,-0.778690), (29465,-0.821366), (29466,-0.999210), (29467,-0.621520), (29468,-0.768707), (29469,-0.818816), (29470,-0.974830), (29471,-0.710476), (29472,-0.883211), (29473,-0.928210), (29474,-1.078650), (29475,-0.535598), (29476,-0.672567), (29477,-0.742650), (29478,-0.908882), (29479,-0.528404), (29480,-0.714609), (29481,-0.751712), (29482,-0.894255), (29483,-0.519815), (29484,-0.677687), (29485,-0.749627), (29486,-0.878235), (29487,-0.620384), (29488,-0.792655), (29489,-0.879922), (29490,-1.039188), (29491,-0.439933), (29492,-0.605236), (29493,-0.666957), (29494,-0.833654), (29495,-0.454570), (29496,-0.748073), (29497,-0.805149), (29498,-0.971846), (29499,-0.540739), (29500,-0.698145), (29501,-0.761259), (29502,-0.914486), (29503,-0.668247), (29504,-0.783850), (29505,-0.844177), (29506,-0.964424), (29507,-0.417657), (29508,-0.604327), (29509,-0.650720), (29510,-0.793263), (29511,-0.452267), (29512,-0.689567), (29513,-0.775442), (29514,-0.927740), (29515,-0.517534), (29516,-0.633601), (29517,-0.715295), (29518,-0.862483), (29519,-0.592554), (29520,-0.729988), (29521,-0.777775), (29522,-0.929143), (29523,-0.429754), (29524,-0.559756), (29525,-0.616368), (29526,-0.796070), (29527,-0.438817), (29528,-0.748114), (29529,-0.802867), (29530,-0.983034), (29531,-0.565397), (29532,-0.703295), (29533,-0.752939), (29534,-0.882476), (29535,-0.648779), (29536,-0.795502), (29537,-0.838643), (29538,-0.999766), (29539,-0.464612), (29540,-0.584394), (29541,-0.665160), (29542,-0.804916), (29543,-0.429548), (29544,-0.730483), (29545,-0.788489), (29546,-0.530173), (29547,-0.498995), (29548,-0.670336), (29549,-0.748314), (29550,-0.908973), (29551,-0.638580), (29552,-0.811780), (29553,-0.866069), (29554,-0.593354), (29555,-0.466026), (29556,-0.662914), (29557,-0.686083), (29558,-0.772886), (29559,-0.495526), (29560,-0.908405), (29561,-0.978022), (29562,-0.725745), (29563,-0.700605), (29564,-0.873805), (29565,-0.907656), (29566,-1.089217), (29567,-0.774698), (29568,-0.912131), (29569,-0.974781), (29570,-1.129401), (29571,-0.577525), (29572,-0.729822), (29573,-0.782253), (29574,-0.951273), (29575,-0.573117), (29576,-0.819707), (29577,-0.873996), (29578,-1.033725), (29579,-0.625842), (29580,-0.771172), (29581,-0.809204), (29582,-0.967075), (29583,-0.698541), (29584,-0.833652), (29585,-0.891657), (29586,-1.098300), (29587,-0.570113), (29588,-0.713120), (29589,-0.771590), (29590,-0.954079), (29591,-0.637702), (29592,-0.855029), (29593,-1.008719), (29594,-1.073227), (29595,-0.830704), (29596,-0.838080), (29597,-0.981087), (29598,-1.028409), (29599,-1.233659), (29600,-0.950725), (29601,-1.091874), (29602,-1.112720), (29603,-0.862765), (29604,-0.687594), (29605,-0.859400), (29606,-0.881175), (29607,-0.950327), (29608,-0.887564), (29609,-1.040326), (29610,-0.712800), (29611,-0.892967), (29612,-0.866434), (29613,-1.028950), (29614,-1.082311), (29615,-1.257368), (29616,-1.006484), (29617,-1.130448), (29618,-0.811748), (29619,-0.924099), (29620,-0.771223), (29621,-0.923056), (29622,-0.892343), (29623,-1.075296), (29624,-0.804904), (29625,-0.939551), (29626,-0.982227), (29627,-0.713228), (29628,-0.721997), (29629,-0.884049), (29630,-0.953202), (29631,-1.166348), (29632,-0.856473), (29633,-1.007842), (29634,-1.067705), (29635,-0.829826), (29636,-0.678344), (29637,-0.839932), (29638,-0.900259), (29639,-0.949439), (29640,-0.725495), (29641,-0.902876), (29642,-0.984570), (29643,-0.714178), (29644,-0.681141), (29645,-0.864096), (29646,-0.905843), (29647,-1.087868), (29648,-0.836984), (29649,-1.019010), (29650,-1.045894), (29651,-0.775501), (29652,-0.616587), (29653,-0.758201), (29654,-0.838037), (29655,-0.896507), (29656,-0.844426), (29657,-1.014375), (29658,-1.056123), (29659,-0.823354), (29660,-0.813543), (29661,-0.982097), (29662,-1.021058), (29663,-1.216089), (29664,-0.921078), (29665,-1.070589), (29666,-1.098866), (29667,-0.885606), (29668,-0.758742), (29669,-0.856229), (29670,-0.942568), (29671,-1.006612), (29672,-0.727859), (29673,-0.893627), (29674,-0.926084), (29675,-0.712824), (29676,-0.687685), (29677,-0.843698), (29678,-0.914245), (29679,-1.092089), (29680,-0.830058), (29681,-0.981426), (29682,-0.979047), (29683,-0.730485), (29684,-0.610589), (29685,-0.795866), (29686,-0.858980), (29687,-0.927204), (29688,-0.681894), (29689,-0.844875), (29690,-0.868043), (29691,-0.633416), (29692,-0.608741), (29693,-0.778689), (29694,-0.843662), (29695,-1.011752), (29696,-0.698626), (29697,-0.880186), (29698,-0.907535), (29699,-0.679411), (29700,-0.510279), (29701,-0.703451), (29702,-0.710362), (29703,-0.818068), (29704,-0.686559), (29705,-0.870907), (29706,-0.919158), (29707,-0.667345), (29708,-0.684474), (29709,-0.839559), (29710,-0.879448), (29711,-1.036390), (29712,-0.775752), (29713,-0.911792), (29714,-0.967940), (29715,-0.670142), (29716,-0.506583), (29717,-0.690466), (29718,-0.745219), (29719,-0.828307), (29720,-0.640595), (29721,-0.715322), (29722,-0.855542), (29723,-0.865240), (29724,-0.608782), (29725,-0.668645), (29726,-0.826516), (29727,-0.547762), (29728,-0.707028), (29729,-0.744595), (29730,-0.876918), (29731,-0.751913), (29732,-0.562807), (29733,-0.592478), (29734,-0.740595), (29735,-0.463235), (29736,-0.792969), (29737,-0.893243), (29738,-1.039967), (29739,-0.588421), (29740,-0.735609), (29741,-0.782931), (29742,-0.964027), (29743,-0.733580), (29744,-0.900742), (29745,-0.943883), (29746,-1.109186), (29747,-0.573567), (29748,-0.703569), (29749,-0.749033), (29750,-0.906440), (29751,-0.554296), (29752,-0.823181), (29753,-0.877006), (29754,-1.015369), (29755,-0.616775), (29756,-0.759319), (29757,-0.803389), (29758,-0.963582), (29759,-0.742427), (29760,-0.891472), (29761,-0.914176), (29762,-1.043713), (29763,-0.546647), (29764,-0.689654), (29765,-0.746730), (29766,-0.887415), (29767,-0.516692), (29768,-0.773965), (29769,-0.822680), (29770,-0.988448), (29771,-0.575920), (29772,-0.731469), (29773,-0.785294), (29774,-0.909722), (29775,-0.656515), (29776,-0.808813), (29777,-0.866353), (29778,-1.010754), (29779,-0.466310), (29780,-0.643690), (29781,-0.676148), (29782,-0.829374), (29783,-0.455864), (29784,-0.592833), (29785,-0.674527), (29786,-0.822644), (29787,-0.791466), (29788,-0.561484), (29789,-0.609270), (29790,-0.778290), (29791,-0.477240), (29792,-0.666698), (29793,-0.744676), (29794,-0.873284), (29795,-0.690681), (29796,-0.471382), (29797,-0.547967), (29798,-0.684937), (29799,-0.447523), (29800,-0.854364), (29801,-0.889608), (29802,-0.664271), (29803,-0.673969), (29804,-0.840201), (29805,-0.890310), (29806,-1.092308), (29807,-0.807981), (29808,-0.971426), (29809,-0.997845), (29810,-0.739994), (29811,-0.587584), (29812,-0.773324), (29813,-0.778377), (29814,-0.896766), (29815,-0.620799), (29816,-0.734080), (29817,-0.816239), (29818,-0.961569), (29819,-0.525351), (29820,-0.676255), (29821,-0.736583), (29822,-0.867513), (29823,-0.634745), (29824,-0.887837), (29825,-0.944913), (29826,-1.089315), (29827,-0.560663), (29828,-0.711567), (29829,-0.779326), (29830,-0.926515), (29831,-0.591557), (29832,-0.722488), (29833,-0.899403), (29834,-0.927216), (29835,-0.663326), (29836,-0.635400), (29837,-0.804419), (29838,-0.858708), (29839,-1.016579), (29840,-0.729930), (29841,-0.876189), (29842,-0.952309), (29843,-0.695386), (29844,-0.528112), (29845,-0.713853), (29846,-0.743524), (29847,-0.851230), (29848,-0.820516), (29849,-0.980246), (29850,-1.016884), (29851,-0.781793), (29852,-0.749221), (29853,-0.926137), (29854,-1.018979), (29855,-1.176386), (29856,-0.899026), (29857,-1.043892), (29858,-1.091677), (29859,-0.853335), (29860,-0.699995), (29861,-0.828603), (29862,-0.889395), (29863,-0.964122), (29864,-0.706735), (29865,-0.851137), (29866,-0.932366), (29867,-0.674515), (29868,-0.686999), (29869,-0.843942), (29870,-0.894515), (29871,-1.091404), (29872,-0.794999), (29873,-0.975166), (29874,-1.028062), (29875,-0.777643), (29876,-0.634986), (29877,-0.790535), (29878,-0.861546), (29879,-0.922338), (29880,-0.796867), (29881,-0.924547), (29882,-0.961649), (29883,-0.741422), (29884,-0.752513), (29885,-0.912707), (29886,-0.943307), (29887,-1.093747), (29888,-0.836824), (29889,-1.012811), (29890,-1.069887), (29891,-0.827364), (29892,-0.678669), (29893,-0.834218), (29894,-0.885720), (29895,-0.962305), (29896,-0.714672), (29897,-0.866505), (29898,-0.903608), (29899,-0.653189), (29900,-0.664744), (29901,-0.841660), (29902,-0.878298), (29903,-1.053356), (29904,-0.781105), (29905,-0.936189), (29906,-1.005807), (29907,-0.755852), (29908,-0.609479), (29909,-0.788717), (29910,-0.818853), (29911,-0.888471), (29912,-0.839642), (29913,-0.991474), (29914,-1.061092), (29915,-0.807886), (29916,-0.790642), (29917,-0.971274), (29918,-1.013951), (29919,-1.188080), (29920,-0.896784), (29921,-1.029109), (29922,-1.077824), (29923,-0.841804), (29924,-0.691251), (29925,-0.851445), (29926,-0.893657), (29927,-0.979531), (29928,-0.709139), (29929,-0.836354), (29930,-0.889714), (29931,-0.675989), (29932,-0.695906), (29933,-0.847274), (29934,-0.850934), (29935,-1.022275), (29936,-0.735161), (29937,-0.896748), (29938,-0.962650), (29939,-0.735455), (29940,-0.559819), (29941,-0.739057), (29942,-0.777554), (29943,-0.824875), (29944,-0.604183), (29945,-0.782028), (29946,-0.835853), (29947,-0.595188), (29948,-0.570048), (29949,-0.758111), (29950,-0.797537), (29951,-0.979098), (29952,-0.678512), (29953,-0.842423), (29954,-0.896247), (29955,-0.648150), (29956,-0.497133), (29957,-0.664294), (29958,-0.717654), (29959,-0.792381), (29960,-0.658085), (29961,-0.851722), (29962,-0.883716), (29963,-0.617504), (29964,-0.622556), (29965,-0.784608), (29966,-0.824962), (29967,-1.007452), (29968,-0.709654), (29969,-0.878209), (29970,-0.949684), (29971,-0.693226), (29972,-0.551963), (29973,-0.718660), (29974,-0.768304), (29975,-0.853250), (29976,-0.657177), (29977,-0.701711), (29978,-0.874446), (29979,-0.872996), (29980,-0.623505), (29981,-0.643887), (29982,-0.846349), (29983,-0.572705), (29984,-0.745905), (29985,-0.783472), (29986,-0.919977), (29987,-0.778249), (29988,-0.526436), (29989,-0.602092), (29990,-0.787369), (29991,-0.442657), (29992,-0.764031), (29993,-0.820177), (29994,-0.968294), (29995,-0.558089), (29996,-0.700167), (29997,-0.776288), (29998,-0.943449), (29999,-0.712074), (30000,-0.835572), (30001,-0.884288), (30002,-1.026831), (30003,-0.475883), (30004,-0.650941), (30005,-0.709411), (30006,-0.859850), (30007,-0.530003), (30008,-0.819790), (30009,-0.830881), (30010,-0.986430), (30011,-0.578547), (30012,-0.758250), (30013,-0.826473), (30014,-0.969017), (30015,-0.696766), (30016,-0.849528), (30017,-0.940512), (30018,-1.089093), (30019,-0.547900), (30020,-0.735964), (30021,-0.783750), (30022,-0.945338), (30023,-0.580652), (30024,-0.823527), (30025,-0.867596), (30026,-1.009675), (30027,-0.576710), (30028,-0.722968), (30029,-0.807449), (30030,-0.939774), (30031,-0.709328), (30032,-0.870915), (30033,-0.881077), (30034,-1.041735), (30035,-0.503793), (30036,-0.634725), (30037,-0.703413), (30038,-0.828769), (30039,-0.478484), (30040,-0.634962), (30041,-0.672065), (30042,-0.815072), (30043,-0.789932), (30044,-0.558093), (30045,-0.639323), (30046,-0.790691), (30047,-0.535627), (30048,-0.686066), (30049,-0.738962), (30050,-0.907981), (30051,-0.762537), (30052,-0.533485), (30053,-0.565478), (30054,-0.688513), (30055,-0.458531), (30056,-0.608041), (30057,-0.758481), (30058,-0.809054), (30059,-0.554918), (30060,-0.569726), (30061,-0.706695), (30062,-0.761913), (30063,-0.975523), (30064,-0.708847), (30065,-0.883440), (30066,-0.922865), (30067,-0.685916), (30068,-0.499597), (30069,-0.664436), (30070,-0.734518), (30071,-0.831540), (30072,-0.794788), (30073,-0.831427), (30074,-0.965609), (30075,-0.580022), (30076,-0.723494), (30077,-0.781498), (30078,-0.937047), (30079,-0.687557), (30080,-0.777612), (30081,-0.966605), (30082,-0.991631), (30083,-0.772797), (30084,-0.597161), (30085,-0.769432), (30086,-0.813038), (30087,-0.876152), (30088,-0.695407), (30089,-0.880683), (30090,-0.919180), (30091,-0.654361), (30092,-0.647337), (30093,-0.804279), (30094,-0.869716), (30095,-1.042916), (30096,-0.764162), (30097,-0.928072), (30098,-0.967962), (30099,-0.712897), (30100,-0.556771), (30101,-0.719287), (30102,-0.762428), (30103,-0.851554), (30104,-0.739090), (30105,-0.867234), (30106,-0.924310), (30107,-0.655310), (30108,-0.675227), (30109,-0.845639), (30110,-0.852086), (30111,-1.039220), (30112,-0.788336), (30113,-0.924841), (30114,-1.002819), (30115,-0.767728), (30116,-0.630181), (30117,-0.802452), (30118,-0.834445), (30119,-0.910101), (30120,-0.989937), (30121,-0.738589), (30122,-0.895531), (30123,-0.543388), (30124,-0.678963), (30125,-0.692376), (30126,-0.853500), (30127,-0.914291), (30128,-1.100961), (30129,-0.831963), (30130,-0.999588), (30131,-0.636761), (30132,-0.800206), (30133,-0.651511), (30134,-0.786622), (30135,-0.759161), (30136,-1.113977), (30137,-0.828721), (30138,-0.943394), (30139,-0.593573), (30140,-0.731936), (30141,-0.728627), (30142,-0.876280), (30143,-0.978412), (30144,-1.130710), (30145,-0.844059), (30146,-0.985673), (30147,-0.639104), (30148,-0.786756), (30149,-0.646422), (30150,-0.810332), (30151,-0.794482), (30152,-0.979759), (30153,-0.703328), (30154,-0.844941), (30155,-0.520668), (30156,-0.665068), (30157,-0.618098), (30158,-0.810806), (30159,-0.871134), (30160,-1.014606), (30161,-0.794843), (30162,-0.924845), (30163,-0.556908), (30164,-0.715709), (30165,-0.586058), (30166,-0.745323), (30167,-0.682559), (30168,-1.126095), (30169,-0.827832), (30170,-0.988955), (30171,-0.600116), (30172,-0.776103), (30173,-0.776047), (30174,-0.926486), (30175,-1.007251), (30176,-1.144220), (30177,-0.887763), (30178,-1.040060), (30179,-0.710212), (30180,-0.848110), (30181,-0.705918), (30182,-0.865183), (30183,-0.816354), (30184,-0.977012), (30185,-0.724271), (30186,-0.851021), (30187,-0.532321), (30188,-0.673470), (30189,-0.639041), (30190,-0.826176), (30191,-0.911121), (30192,-1.069922), (30193,-0.774446), (30194,-0.910021), (30195,-0.567632), (30196,-0.736652), (30197,-0.607930), (30198,-0.759298), (30199,-0.725798), (30200,-0.949627), (30201,-0.670409), (30202,-0.779509), (30203,-0.481711), (30204,-0.631221), (30205,-0.619088), (30206,-0.770921), (30207,-0.824281), (30208,-0.966360), (30209,-0.706185), (30210,-0.848729), (30211,-0.518881), (30212,-0.672572), (30213,-0.521089), (30214,-0.680355), (30215,-0.649177), (30216,-0.957544), (30217,-0.673217), (30218,-0.839914), (30219,-0.484054), (30220,-0.615449), (30221,-0.652087), (30222,-0.758864), (30223,-0.845203), (30224,-0.984030), (30225,-0.718283), (30226,-0.913778), (30227,-0.565351), (30228,-0.709287), (30229,-0.527148), (30230,-0.705457), (30231,-0.684963), (30232,-0.506540), (30233,-0.650477), (30234,-0.708946), (30235,-0.847309), (30236,-0.438961), (30237,-0.608445), (30238,-0.641367), (30239,-0.805277), (30240,-0.569257), (30241,-0.687647), (30242,-0.752154), (30243,-0.909097), (30244,-0.367904), (30245,-0.487222), (30246,-0.555911), (30247,-0.711924), (30248,-0.614323), (30249,-0.804709), (30250,-0.808369), (30251,-0.590928), (30252,-0.596910), (30253,-0.732950), (30254,-0.810928), (30255,-0.968799), (30256,-0.694691), (30257,-0.853027), (30258,-0.914748), (30259,-0.651323), (30260,-0.491479), (30261,-0.648887), (30262,-0.695744), (30263,-0.795553), (30264,-0.597622), (30265,-0.774537), (30266,-0.843226), (30267,-0.583981), (30268,-0.571383), (30269,-0.728325), (30270,-0.772860), (30271,-0.933054), (30272,-0.650584), (30273,-0.799166), (30274,-0.867854), (30275,-0.650414), (30276,-0.487319), (30277,-0.656338), (30278,-0.688797), (30279,-0.735189), (30280,-0.572095), (30281,-0.733218), (30282,-0.813054), (30283,-0.590504), (30284,-0.571403), (30285,-0.752035), (30286,-0.758945), (30287,-0.911707), (30288,-0.650605), (30289,-0.798722), (30290,-0.858120), (30291,-0.596553), (30292,-0.443213), (30293,-0.613625), (30294,-0.682778), (30295,-0.711985), (30296,-0.420690), (30297,-0.557194), (30298,-0.607767), (30299,-0.741485), (30300,-0.346143), (30301,-0.528633), (30302,-0.588496), (30303,-0.731968), (30304,-0.468078), (30305,-0.640349), (30306,-0.675594), (30307,-0.868767), (30308,-0.299240), (30309,-0.434816), (30310,-0.527658), (30311,-0.694354), (30312,-0.539156), (30313,-0.676590), (30314,-0.719731), (30315,-0.491607), (30316,-0.466003), (30317,-0.606688), (30318,-0.690241), (30319,-0.831390), (30320,-0.547992), (30321,-0.751848), (30322,-0.797312), (30323,-0.552466), (30324,-0.413525), (30325,-0.575578), (30326,-0.619183), (30327,-0.713419), (30328,-0.585161), (30329,-0.744891), (30330,-0.789890), (30331,-0.545974), (30332,-0.541736), (30333,-0.668022), (30334,-0.723705), (30335,-0.874144), (30336,-0.790943), (30337,-0.955782), (30338,-1.004961), (30339,-0.783805), (30340,-0.633716), (30341,-0.778582), (30342,-0.822652), (30343,-0.929893), (30344,-0.746361), (30345,-0.899588), (30346,-0.936690), (30347,-0.697884), (30348,-0.669028), (30349,-0.825506), (30350,-0.890478), (30351,-1.079006), (30352,-0.807685), (30353,-0.963698), (30354,-1.009162), (30355,-0.780109), (30356,-0.637453), (30357,-0.805078), (30358,-0.870980), (30359,-0.945707), (30360,-1.189045), (30361,-0.884744), (30362,-1.019391), (30363,-0.686756), (30364,-0.851594), (30365,-0.826920), (30366,-0.991759), (30367,-1.056267), (30368,-1.214602), (30369,-0.916805), (30370,-1.037981), (30371,-0.711385), (30372,-0.891087), (30373,-0.732173), (30374,-0.880755), (30375,-0.837035), (30376,-1.046930), (30377,-0.772357), (30378,-0.928835), (30379,-0.592019), (30380,-0.759645), (30381,-0.735899), (30382,-0.866830), (30383,-0.931338), (30384,-1.082242), (30385,-0.834145), (30386,-0.992945), (30387,-0.637085), (30388,-0.795421), (30389,-0.656481), (30390,-0.794843), (30391,-0.768775), (30392,-1.092006), (30393,-0.798853), (30394,-0.943254), (30395,-0.623626), (30396,-0.742944), (30397,-0.763789), (30398,-0.946743), (30399,-1.018683), (30400,-1.136608), (30401,-0.893620), (30402,-1.022228), (30403,-0.714676), (30404,-0.874406), (30405,-0.732213), (30406,-0.878937), (30407,-0.827322), (30408,-1.018637), (30409,-0.748708), (30410,-0.901006), (30411,-0.537714), (30412,-0.658426), (30413,-0.701567), (30414,-0.866406), (30415,-0.915121), (30416,-1.073921), (30417,-0.825824), (30418,-0.967438), (30419,-0.617617), (30420,-0.734613), (30421,-0.591957), (30422,-0.773052), (30423,-0.741410), (30424,-1.175656), (30425,-0.879716), (30426,-1.076140), (30427,-0.728177), (30428,-0.836347), (30429,-0.782410), (30430,-0.977440), (30431,-1.032658), (30432,-1.171021), (30433,-0.868114), (30434,-1.022269), (30435,-0.718897), (30436,-0.848899), (30437,-0.702527), (30438,-0.825561), (30439,-0.828291), (30440,-0.956899), (30441,-0.715770), (30442,-0.855061), (30443,-0.515923), (30444,-0.673795), (30445,-0.705788), (30446,-0.836719), (30447,-0.896117), (30448,-1.087432), (30449,-0.791492), (30450,-0.960047), (30451,-0.645527), (30452,-0.783426), (30453,-0.610577), (30454,-0.758229), (30455,-0.765140), (30456,-0.831041), (30457,-0.573655), (30458,-0.746855), (30459,-0.805788), (30460,-0.553975), (30461,-0.496321), (30462,-0.632361), (30463,-0.704301), (30464,-0.869605), (30465,-0.588993), (30466,-0.736181), (30467,-0.800225), (30468,-0.514039), (30469,-0.365809), (30470,-0.514855), (30471,-0.558460), (30472,-0.768355), (30473,-0.491459), (30474,-0.650260), (30475,-0.697581), (30476,-0.484786), (30477,-0.441531), (30478,-0.634240), (30479,-0.685277), (30480,-0.866373), (30481,-0.584369), (30482,-0.777541), (30483,-0.840656), (30484,-0.571657), (30485,-0.414136), (30486,-0.579904), (30487,-0.615148), (30488,-0.500362), (30489,-0.632686), (30490,-0.654461), (30491,-0.805365), (30492,-0.425351), (30493,-0.615273), (30494,-0.673278), (30495,-0.820930), (30496,-0.539389), (30497,-0.681003), (30498,-0.734828), (30499,-0.907099), (30500,-0.371944), (30501,-0.518668), (30502,-0.577602), (30503,-0.707604), (30504,-0.604894), (30505,-0.773913), (30506,-0.832382), (30507,-0.582892), (30508,-0.570294), (30509,-0.717946), (30510,-0.772235), (30511,-0.954260), (30512,-0.674578), (30513,-0.841274), (30514,-0.889525), (30515,-0.673943), (30516,-0.478798), (30517,-0.656643), (30518,-0.691888), (30519,-0.768937), (30520,-0.464172), (30521,-0.606715), (30522,-0.676332), (30523,-0.796115), (30524,-0.383123), (30525,-0.547961), (30526,-0.633836), (30527,-0.757799), (30528,-0.504593), (30529,-0.662000), (30530,-0.691670), (30531,-0.867658), (30532,-0.297201), (30533,-0.443925), (30534,-0.514936), (30535,-0.678845), (30536,-0.379190), (30537,-0.547280), (30538,-0.617826), (30539,-0.748757), (30540,-0.354808), (30541,-0.539156), (30542,-0.578582), (30543,-0.748995), (30544,-0.499504), (30545,-0.667130), (30546,-0.708413), (30547,-0.846775), (30548,-0.312550), (30549,-0.452771), (30550,-0.515885), (30551,-0.687227), (30552,-0.403363), (30553,-0.542191), (30554,-0.589512), (30555,-0.735771), (30556,-0.358081), (30557,-0.497372), (30558,-0.585105), (30559,-0.750408), (30560,-0.512065), (30561,-0.661576), (30562,-0.695428), (30563,-0.889065), (30564,-0.361807), (30565,-0.503421), (30566,-0.592082), (30567,-0.726729), (30568,-0.560847), (30569,-0.759130), (30570,-0.797161), (30571,-0.532808), (30572,-0.521603), (30573,-0.695732), (30574,-0.722151), (30575,-0.905105), (30576,-0.626351), (30577,-0.793977), (30578,-0.801817), (30579,-0.544430), (30580,-0.396664), (30581,-0.560109), (30582,-0.624153), (30583,-0.680764), (30584,-0.560403), (30585,-0.710843), (30586,-0.765132), (30587,-0.549085), (30588,-0.525339), (30589,-0.693894), (30590,-0.776053), (30591,-0.953897), (30592,-0.877663), (30593,-1.037392), (30594,-1.096791), (30595,-0.840798), (30596,-0.689780), (30597,-0.843006), (30598,-0.872678), (30599,-0.968771), (30600,-0.802890), (30601,-0.909667), (30602,-0.978820), (30603,-0.727936), (30604,-0.699080), (30605,-0.870422), (30606,-0.946078), (30607,-1.134606), (30608,-0.832628), (30609,-0.996537), (30610,-1.036427), (30611,-0.792046), (30612,-0.646138), (30613,-0.817945), (30614,-0.875020), (30615,-0.942316), (30616,-0.958516), (30617,-0.648641), (30618,-0.802797), (30619,-0.885420), (30620,-0.648471), (30621,-0.642375), (30622,-0.789099), (30623,-0.859181), (30624,-1.004511), (30625,-0.706248), (30626,-0.889667), (30627,-0.910977), (30628,-0.687498), (30629,-0.529513), (30630,-0.701784), (30631,-0.739351), (30632,-0.988264), (30633,-0.709510), (30634,-0.841834), (30635,-0.512916), (30636,-0.663819), (30637,-0.684665), (30638,-0.819776), (30639,-0.916334), (30640,-1.066309), (30641,-0.754576), (30642,-0.930563), (30643,-0.619759), (30644,-0.765554), (30645,-0.639619), (30646,-0.785878), (30647,-0.735191), (30648,-1.137851), (30649,-0.855846), (30650,-1.003963), (30651,-0.682012), (30652,-0.820839), (30653,-0.811028), (30654,-0.985156), (30655,-1.073353), (30656,-1.211251), (30657,-0.961297), (30658,-1.067609), (30659,-0.718252), (30660,-0.883556), (30661,-0.719997), (30662,-0.871365), (30663,-0.843903), (30664,-1.032896), (30665,-0.781547), (30666,-0.903653), (30667,-0.554761), (30668,-0.718670), (30669,-0.702356), (30670,-0.876020), (30671,-0.940528), (30672,-1.099329), (30673,-0.796421), (30674,-0.971479), (30675,-0.639309), (30676,-0.784639), (30677,-0.636873), (30678,-0.835620), (30679,-0.793293), (30680,-0.985073), (30681,-0.723041), (30682,-0.880448), (30683,-0.924983), (30684,-0.688963), (30685,-0.682403), (30686,-0.833772), (30687,-0.854617), (30688,-1.049648), (30689,-0.773217), (30690,-0.881388), (30691,-0.931960), (30692,-0.693153), (30693,-0.511015), (30694,-0.693040), (30695,-0.771018), (30696,-0.852712), (30697,-0.564669), (30698,-0.729508), (30699,-0.785655), (30700,-0.561711), (30701,-0.512883), (30702,-0.667967), (30703,-0.721792), (30704,-0.908926), (30705,-0.616238), (30706,-0.777826), (30707,-0.825147), (30708,-0.598881), (30709,-0.416742), (30710,-0.579723), (30711,-0.620542), (30712,-0.754260), (30713,-0.481080), (30714,-0.629197), (30715,-0.657010), (30716,-0.410771), (30717,-0.409321), (30718,-0.586701), (30719,-0.649351), (30720,-1.125865), (30721,-1.250758), (30722,-0.982223), (30723,-0.769428), (30724,-0.825575), (30725,-0.987627), (30726,-0.786444), (30727,-0.867674), (30728,-1.127269), (30729,-1.289321), (30730,-1.014283), (30731,-0.741104), (30732,-0.822798), (30733,-0.987637), (30734,-0.978290), (30735,-1.151954), (30736,-1.231791), (30737,-1.383159), (30738,-1.088148), (30739,-0.843767), (30740,-0.876690), (30741,-1.070792), (30742,-0.896550), (30743,-0.967560), (30744,-1.200680), (30745,-0.946080), (30746,-1.096520), (30747,-0.729512), (30748,-0.889241), (30749,-0.866888), (30750,-1.020579), (30751,-1.085087), (30752,-1.242030), (30753,-0.971173), (30754,-1.112323), (30755,-0.783403), (30756,-0.900399), (30757,-0.777716), (30758,-0.915150), (30759,-0.900694), (30760,-1.081789), (30761,-0.805358), (30762,-0.987848), (30763,-0.638491), (30764,-0.801937), (30765,-0.813492), (30766,-0.946281), (30767,-1.015434), (30768,-1.180272), (30769,-0.910809), (30770,-1.027340), (30771,-0.696563), (30772,-0.848396), (30773,-0.688088), (30774,-0.839922), (30775,-0.817569), (30776,-1.146839), (30777,-0.888523), (30778,-1.023634), (30779,-0.687283), (30780,-0.825646), (30781,-0.831163), (30782,-0.986247), (30783,-1.068406), (30784,-1.198408), (30785,-0.971213), (30786,-1.122117), (30787,-0.807133), (30788,-0.950605), (30789,-0.809342), (30790,-0.940737), (30791,-0.912346), (30792,-1.189128), (30793,-0.901085), (30794,-1.049202), (30795,-0.695200), (30796,-0.859110), (30797,-0.852550), (30798,-0.989983), (30799,-1.060995), (30800,-1.177061), (30801,-0.940577), (30802,-1.091946), (30803,-0.738408), (30804,-0.884203), (30805,-0.779170), (30806,-0.899882), (30807,-0.869168), (30808,-1.117616), (30809,-0.842114), (30810,-0.975368), (30811,-0.662706), (30812,-0.778308), (30813,-0.790328), (30814,-0.952380), (30815,-1.028500), (30816,-1.171044), (30817,-0.905295), (30818,-1.057593), (30819,-0.685011), (30820,-0.823839), (30821,-0.671892), (30822,-0.819080), (30823,-0.841784), (30824,-1.217039), (30825,-0.922492), (30826,-0.676717), (30827,-0.773276), (30828,-0.954372), (30829,-0.919478), (30830,-1.088962), (30831,-1.133032), (30832,-1.310412), (30833,-1.037232), (30834,-0.818399), (30835,-0.863863), (30836,-0.988754), (30837,-0.833092), (30838,-0.934760), (30839,-0.968147), (30840,-1.177577), (30841,-0.869096), (30842,-1.025109), (30843,-0.724989), (30844,-0.869854), (30845,-0.842857), (30846,-0.990045), (30847,-1.053623), (30848,-1.396364), (30849,-1.122255), (30850,-0.907602), (30851,-0.949814), (30852,-1.112330), (30853,-0.965494), (30854,-1.037897), (30855,-1.063853), (30856,-1.206860), (30857,-1.352655), (30858,-0.686977), (30859,-0.824875), (30860,-0.897744), (30861,-1.068621), (30862,-1.081571), (30863,-1.184631), (30864,-1.231024), (30865,-1.421410), (30866,-0.759448), (30867,-0.895024), (30868,-0.925160), (30869,-1.085354), (30870,-0.841901), (30871,-0.996521), (30872,-1.251472), (30873,-1.413524), (30874,-0.772000), (30875,-0.947522), (30876,-0.986483), (30877,-1.162470), (30878,-1.169845), (30879,-1.325393), (30880,-1.369928), (30881,-1.541270), (30882,-0.875592), (30883,-1.008845), (30884,-1.051058), (30885,-1.181059), (30886,-0.979412), (30887,-1.103375), (30888,-1.156271), (30889,-1.344334), (30890,-0.687947), (30891,-0.819342), (30892,-0.903823), (30893,-1.047760), (30894,-1.056528), (30895,-1.223690), (30896,-1.303525), (30897,-1.491125), (30898,-0.781320), (30899,-0.938263), (30900,-1.005093), (30901,-1.126269), (30902,-0.911616), (30903,-1.071345), (30904,-1.306323), (30905,-1.470697), (30906,-0.738132), (30907,-0.901578), (30908,-0.957725), (30909,-1.139285), (30910,-1.143873), (30911,-1.325434), (30912,-1.362072), (30913,-1.507867), (30914,-0.819429), (30915,-0.953146), (30916,-0.991643), (30917,-1.128147), (30918,-0.915352), (30919,-1.049999), (30920,-1.147951), (30921,-1.276559), (30922,-0.620171), (30923,-0.748779), (30924,-0.861595), (30925,-1.036188), (30926,-1.023125), (30927,-1.194002), (30928,-1.257117), (30929,-1.388512), (30930,-0.701003), (30931,-0.881635), (30932,-0.940569), (30933,-1.102156), (30934,-0.865207), (30935,-0.999389), (30936,-1.291964), (30937,-1.460984), (30938,-0.777190), (30939,-0.917875), (30940,-0.997712), (30941,-1.146758), (30942,-1.144379), (30943,-1.285528), (30944,-1.322166), (30945,-1.516733), (30946,-0.829689), (30947,-0.974089), (30948,-1.042778), (30949,-1.189037), (30950,-0.982280), (30951,-1.128075), (30952,-1.169358), (30953,-1.357886), (30954,-0.698711), (30955,-0.829642), (30956,-0.895079), (30957,-1.073852), (30958,-1.069151), (30959,-1.213551), (30960,-1.311039), (30961,-1.461014), (30962,-0.774899), (30963,-0.929518), (30964,-1.020038), (30965,-1.142143), (30966,-0.882434), (30967,-1.044486), (30968,-1.138257), (30969,-1.313315), (30970,-0.648566), (30971,-0.748376), (30972,-0.804987), (30973,-0.993515), (30974,-0.996710), (30975,-1.141575), (30976,-1.226986), (30977,-1.367671), (30978,-0.702458), (30979,-0.845001), (30980,-0.895109), (30981,-1.075277), (30982,-0.855513), (30983,-0.980870), (30984,-1.185191), (30985,-1.335631), (30986,-0.651373), (30987,-0.818999), (30988,-0.847741), (30989,-1.007935), (30990,-1.047825), (30991,-1.168536), (30992,-1.239547), (30993,-1.396025), (30994,-0.728954), (30995,-0.876142), (30996,-0.921141), (30997,-1.072045), (30998,-0.852747), (30999,-1.011547), (31000,-1.154555), (31001,-0.870227), (31002,-1.024382), (31003,-0.718688), (31004,-0.877953), (31005,-0.901121), (31006,-1.059457), (31007,-1.128610), (31008,-1.293449), (31009,-1.008193), (31010,-1.143768), (31011,-0.825068), (31012,-0.919304), (31013,-0.759925), (31014,-0.934518), (31015,-0.891263), (31016,-1.307858), (31017,-1.026782), (31018,-0.766609), (31019,-0.799995), (31020,-0.981091), (31021,-0.981035), (31022,-1.166311), (31023,-1.223852), (31024,-1.405413), (31025,-1.128052), (31026,-0.896677), (31027,-0.937496), (31028,-1.076323), (31029,-0.922054), (31030,-0.998639), (31031,-1.054786), (31032,-1.283725), (31033,-1.007294), (31034,-0.769881), (31035,-0.824634), (31036,-0.964390), (31037,-0.939251), (31038,-1.121740), (31039,-1.203434), (31040,-1.364093), (31041,-1.069546), (31042,-0.814946), (31043,-0.865055), (31044,-1.017817), (31045,-0.826853), (31046,-0.902973), (31047,-0.934038), (31048,-1.209426), (31049,-0.931602), (31050,-0.714161), (31051,-0.782850), (31052,-0.950011), (31053,-0.954134), (31054,-1.130122), (31055,-1.156540), (31056,-1.292116), (31057,-1.023117), (31058,-0.787097), (31059,-0.846496), (31060,-1.009941), (31061,-0.866355), (31062,-0.918322), (31063,-0.983294), (31064,-1.082640), (31065,-0.819214), (31066,-0.941784), (31067,-0.626800), (31068,-0.756337), (31069,-0.751635), (31070,-0.880708), (31071,-0.984233), (31072,-1.137924), (31073,-0.876357), (31074,-1.032370), (31075,-0.702523), (31076,-0.894302), (31077,-0.708912), (31078,-0.831482), (31079,-0.808665), (31080,-1.163482), (31081,-0.899592), (31082,-0.664965), (31083,-0.707177), (31084,-0.865978), (31085,-0.822259), (31086,-0.983846), (31087,-1.014446), (31088,-1.185788), (31089,-0.869875), (31090,-0.628281), (31091,-0.693717), (31092,-0.854840), (31093,-0.717757), (31094,-0.818496), (31095,-0.874643), (31096,-1.214596), (31097,-0.921444), (31098,-0.672882), (31099,-0.740177), (31100,-0.893403), (31101,-0.888702), (31102,-1.070262), (31103,-1.105507), (31104,-1.385540), (31105,-1.107251), (31106,-0.874947), (31107,-0.945958), (31108,-1.110797), (31109,-0.974179), (31110,-1.038222), (31111,-1.086009), (31112,-1.350713), (31113,-1.072889), (31114,-0.900969), (31115,-0.926459), (31116,-1.072254), (31117,-1.068946), (31118,-1.245862), (31119,-1.311298), (31120,-1.446874), (31121,-1.180662), (31122,-0.939068), (31123,-0.953875), (31124,-1.091309), (31125,-0.962586), (31126,-1.035456), (31127,-1.071165), (31128,-1.289421), (31129,-1.426389), (31130,-0.761176), (31131,-0.956208), (31132,-0.995168), (31133,-1.155827), (31134,-1.159950), (31135,-1.312712), (31136,-1.360498), (31137,-1.514654), (31138,-0.851299), (31139,-1.021712), (31140,-1.058349), (31141,-1.179526), (31142,-0.984846), (31143,-1.145504), (31144,-1.253210), (31145,-1.392966), (31146,-0.707780), (31147,-0.865651), (31148,-0.949203), (31149,-1.080135), (31150,-1.083329), (31151,-1.250025), (31152,-1.297348), (31153,-1.464044), (31154,-0.790470), (31155,-0.940909), (31156,-1.012385), (31157,-1.166540), (31158,-0.915192), (31159,-1.056342), (31160,-1.265307), (31161,-1.397632), (31162,-0.723593), (31163,-0.877748), (31164,-0.940863), (31165,-1.096876), (31166,-1.120045), (31167,-1.293708), (31168,-1.333133), (31169,-1.489147), (31170,-0.828579), (31171,-0.982270), (31172,-0.992896), (31173,-1.170741), (31174,-0.918928), (31175,-1.055898), (31176,-1.184970), (31177,-1.353989), (31178,-0.667410), (31179,-0.820636), (31180,-0.888395), (31181,-1.037441), (31182,-1.051319), (31183,-1.239847), (31184,-1.263016), (31185,-1.379547), (31186,-0.725017), (31187,-0.894037), (31188,-0.969692), (31189,-1.117809), (31190,-0.884112), (31191,-0.998321), (31192,-1.341060), (31193,-1.490571), (31194,-0.795630), (31195,-0.931206), (31196,-0.977599), (31197,-1.165198), (31198,-1.172109), (31199,-1.346702), (31200,-1.343393), (31201,-1.487794), (31202,-0.840697), (31203,-1.025044), (31204,-1.065863), (31205,-1.209799), (31206,-0.981211), (31207,-1.136296), (31208,-1.205913), (31209,-1.355423), (31210,-0.693462), (31211,-0.852262), (31212,-0.913054), (31213,-1.041662), (31214,-1.049038), (31215,-1.212018), (31216,-1.281636), (31217,-1.438114), (31218,-0.802164), (31219,-0.939133), (31220,-0.991100), (31221,-1.139681), (31222,-0.907841), (31223,-1.043417), (31224,-1.172954), (31225,-1.322000), (31226,-0.648890), (31227,-0.794220), (31228,-0.884741), (31229,-1.046328), (31230,-1.035123), (31231,-1.161873), (31232,-1.196189), (31233,-1.364744), (31234,-0.671196), (31235,-0.790979), (31236,-0.873603), (31237,-1.004069), (31238,-0.768049), (31239,-0.938461), (31240,-1.192018), (31241,-1.358251), (31242,-0.641943), (31243,-0.777519), (31244,-0.840169), (31245,-0.994325), (31246,-1.024460), (31247,-1.185582), (31248,-1.269135), (31249,-1.417716), (31250,-0.726027), (31251,-0.864854), (31252,-0.907531), (31253,-1.060757), (31254,-0.815912), (31255,-0.975177), (31256,-1.108895), (31257,-0.850114), (31258,-0.994051), (31259,-0.635868), (31260,-0.832757), (31261,-0.821088), (31262,-0.946909), (31263,-1.031391), (31264,-1.235247), (31265,-0.917940), (31266,-1.072096), (31267,-0.727384), (31268,-0.857386), (31269,-0.703581), (31270,-0.842408), (31271,-0.838171), (31272,-1.272881), (31273,-0.977870), (31274,-0.734883), (31275,-0.811933), (31276,-0.989312), (31277,-0.981359), (31278,-1.147127), (31279,-1.194448), (31280,-1.343030), (31281,-1.081927), (31282,-0.838475), (31283,-0.887655), (31284,-1.049243), (31285,-0.874536), (31286,-0.962733), (31287,-1.005410), (31288,-1.291481), (31289,-1.006225), (31290,-0.755806), (31291,-0.828210), (31292,-0.979578), (31293,-0.945613), (31294,-1.105807), (31295,-1.164741), (31296,-1.331903), (31297,-1.038285), (31298,-0.831064), (31299,-0.905326), (31300,-1.067378), (31301,-0.918218), (31302,-0.981333), (31303,-1.035157), (31304,-1.280354), (31305,-0.982556), (31306,-0.751181), (31307,-0.801754), (31308,-0.973560), (31309,-0.967929), (31310,-1.131839), (31311,-1.201921), (31312,-1.359328), (31313,-1.059672), (31314,-0.832942), (31315,-0.839388), (31316,-1.019555), (31317,-0.869467), (31318,-0.962309), (31319,-1.000805), (31320,-1.094576), (31321,-0.830222), (31322,-1.007138), (31323,-0.669393), (31324,-0.847702), (31325,-0.817454), (31326,-0.977183), (31327,-1.049123), (31328,-1.208852), (31329,-0.918486), (31330,-1.084254), (31331,-0.731181), (31332,-0.865363), (31333,-0.725958), (31334,-0.869895), (31335,-0.833143), (31336,-1.210720), (31337,-0.922677), (31338,-0.701520), (31339,-0.726547), (31340,-0.916468), (31341,-0.886684), (31342,-1.091004), (31343,-1.118817), (31344,-1.258109), (31345,-0.978891), (31346,-0.747515), (31347,-0.841287), (31348,-0.997765), (31349,-0.829096), (31350,-0.894069), (31351,-0.962757), (31352,-1.297136), (31353,-1.022563), (31354,-0.755422), (31355,-0.804602), (31356,-0.960615), (31357,-0.948017), (31358,-1.163486), (31359,-1.199195), (31360,-1.334306), (31361,-1.459198), (31362,-0.771225), (31363,-0.927703), (31364,-1.029370), (31365,-1.177952), (31366,-0.934500), (31367,-1.110951), (31368,-1.419783), (31369,-1.176796), (31370,-0.884572), (31371,-1.028508), (31372,-1.081869), (31373,-1.275506), (31374,-1.223426), (31375,-1.381297), (31376,-1.436980), (31377,-1.209320), (31378,-0.925458), (31379,-1.061498), (31380,-1.100923), (31381,-1.217919), (31382,-1.038567), (31383,-1.208051), (31384,-1.266520), (31385,-1.438327), (31386,-0.762430), (31387,-0.917050), (31388,-0.970875), (31389,-1.115276), (31390,-1.118470), (31391,-1.280522), (31392,-1.372435), (31393,-1.514514), (31394,-0.885996), (31395,-1.042474), (31396,-1.115343), (31397,-1.186818), (31398,-0.948476), (31399,-1.106811), (31400,-1.389167), (31401,-1.068144), (31402,-1.230197), (31403,-0.960268), (31404,-1.106527), (31405,-1.188686), (31406,-1.344235), (31407,-1.324205), (31408,-1.483934), (31409,-1.142939), (31410,-1.283159), (31411,-0.995115), (31412,-1.127440), (31413,-1.105087), (31414,-1.256920), (31415,-1.136559), (31416,-1.328803), (31417,-1.481101), (31418,-0.789876), (31419,-0.965398), (31420,-1.021081), (31421,-1.181275), (31422,-1.209087), (31423,-1.337231), (31424,-1.367367), (31425,-1.523844), (31426,-0.834942), (31427,-1.003497), (31428,-1.086585), (31429,-1.216586), (31430,-0.974063), (31431,-1.128683), (31432,-1.369699), (31433,-0.989221), (31434,-1.151273), (31435,-0.870662), (31436,-1.045255), (31437,-1.140884), (31438,-1.284355), (31439,-1.266184), (31440,-1.456105), (31441,-1.087240), (31442,-1.226996), (31443,-0.947778), (31444,-1.097753), (31445,-1.089335), (31446,-1.278792), (31447,-1.110588), (31448,-1.247557), (31449,-1.402641), (31450,-0.734177), (31451,-0.839096), (31452,-0.892456), (31453,-1.069836), (31454,-1.093004), (31455,-1.231831), (31456,-1.297733), (31457,-1.443992), (31458,-0.770883), (31459,-0.922251), (31460,-0.989546), (31461,-1.158565), (31462,-0.938337), (31463,-1.086454), (31464,-1.117983), (31465,-1.155551), (31466,-0.909776), (31467,-0.611050), (31468,-0.769386), (31469,-0.812062), (31470,-0.997339), (31471,-0.972199), (31472,-1.121245), (31473,-1.165780), (31474,-0.911180), (31475,-0.647755), (31476,-0.836747), (31477,-0.865025), (31478,-0.943003), (31479,-0.756684), (31480,-0.996771), (31481,-1.123057), (31482,-0.450412), (31483,-0.626863), (31484,-0.695086), (31485,-0.865964), (31486,-0.880306), (31487,-1.037249), (31488,-1.041372), (31489,-1.208998), (31490,-0.546572), (31491,-0.700263), (31492,-0.752694), (31493,-0.902204), (31494,-0.696377), (31495,-0.864932), (31496,-1.078542), (31497,-1.122148), (31498,-0.858723), (31499,-0.586472), (31500,-0.771748), (31501,-0.828360), (31502,-1.019211), (31503,-1.016367), (31504,-1.178419), (31505,-1.191832), (31506,-1.006442), (31507,-0.678452), (31508,-0.838646), (31509,-0.859027), (31510,-0.919354), (31511,-0.757189), (31512,-1.174713), (31513,-1.313540), (31514,-0.643682), (31515,-0.779257), (31516,-0.856772), (31517,-0.997921), (31518,-1.039204), (31519,-1.220764), (31520,-1.249042), (31521,-1.403662), (31522,-0.731481), (31523,-0.870773), (31524,-0.902302), (31525,-1.042522), (31526,-0.797677), (31527,-0.963909), (31528,-1.033062), (31529,-1.197436), (31530,-0.503889), (31531,-0.679876), (31532,-0.729056), (31533,-0.885533), (31534,-0.893373), (31535,-1.065644), (31536,-1.095779), (31537,-1.264799), (31538,-0.581005), (31539,-0.768605), (31540,-0.839615), (31541,-1.003061), (31542,-0.740100), (31543,-0.857560), (31544,-1.074423), (31545,-1.223468), (31546,-0.574049), (31547,-0.690580), (31548,-0.761590), (31549,-0.921784), (31550,-0.951919), (31551,-1.074954), (31552,-1.118095), (31553,-1.273644), (31554,-0.568949), (31555,-0.775592), (31556,-0.806657), (31557,-0.954774), (31558,-0.700638), (31559,-0.885450), (31560,-1.048431), (31561,-1.223489), (31562,-0.558740), (31563,-0.685491), (31564,-0.730025), (31565,-0.883252), (31566,-0.896665), (31567,-1.061504), (31568,-1.140876), (31569,-1.288993), (31570,-0.591265), (31571,-0.731486), (31572,-0.799245), (31573,-0.995205), (31574,-0.741070), (31575,-0.897547), (31576,-1.185477), (31577,-1.319195), (31578,-0.682781), (31579,-0.819285), (31580,-0.881935), (31581,-1.024014), (31582,-1.049504), (31583,-1.196228), (31584,-1.279315), (31585,-1.386557), (31586,-0.709267), (31587,-0.857848), (31588,-0.945116), (31589,-1.081621), (31590,-0.835382), (31591,-0.958417), (31592,-1.211045), (31593,-1.005217), (31594,-0.691162), (31595,-0.869006), (31596,-0.902393), (31597,-1.086741), (31598,-1.061137), (31599,-1.198570), (31600,-1.279800), (31601,-1.062824), (31602,-0.782213), (31603,-0.922898), (31604,-0.970220), (31605,-1.016612), (31606,-0.866524), (31607,-1.055516), (31608,-1.123740), (31609,-1.296011), (31610,-0.627546), (31611,-0.774734), (31612,-0.835527), (31613,-0.968315), (31614,-1.006347), (31615,-1.136813), (31616,-1.423349), (31617,-1.587724), (31618,-0.889067), (31619,-1.071092), (31620,-1.100298), (31621,-1.246557), (31622,-1.006821), (31623,-1.204175), (31624,-1.238955), (31625,-1.290457), (31626,-1.050721), (31627,-0.783115), (31628,-0.947954), (31629,-1.000850), (31630,-1.198203), (31631,-1.167025), (31632,-1.321645), (31633,-1.383831), (31634,-1.145488), (31635,-0.863483), (31636,-0.996736), (31637,-1.051490), (31638,-1.115069), (31639,-0.963587), (31640,-1.367640), (31641,-1.407994), (31642,-1.134351), (31643,-0.889970), (31644,-1.030655), (31645,-1.058467), (31646,-1.258143), (31647,-1.247868), (31648,-1.412707), (31649,-1.472105), (31650,-1.219363), (31651,-0.970802), (31652,-1.144930), (31653,-1.178317), (31654,-1.233535), (31655,-1.058364), (31656,-1.295664), (31657,-1.338805), (31658,-1.083741), (31659,-0.829606), (31660,-0.988406), (31661,-1.011573), (31662,-1.222397), (31663,-1.201903), (31664,-1.345840), (31665,-1.391303), (31666,-1.142277), (31667,-0.879781), (31668,-1.010711), (31669,-1.052460), (31670,-1.100246), (31671,-0.952479), (31672,-1.406234), (31673,-1.441479), (31674,-1.211032), (31675,-0.906732), (31676,-1.063210), (31677,-1.122608), (31678,-1.313459), (31679,-1.304577), (31680,-1.491247), (31681,-1.533923), (31682,-1.305335), (31683,-1.009860), (31684,-1.171912), (31685,-1.203441), (31686,-1.288851), (31687,-1.123434), (31688,-1.252042), (31689,-1.309118), (31690,-1.067059), (31691,-0.771584), (31692,-0.963363), (31693,-0.998144), (31694,-1.154157), (31695,-1.121121), (31696,-1.292463), (31697,-1.308664), (31698,-1.064747), (31699,-0.772988), (31700,-0.948510), (31701,-0.983290), (31702,-1.094248), (31703,-0.905606), (31704,-1.344032), (31705,-1.372310), (31706,-1.125142), (31707,-0.832918), (31708,-1.012156), (31709,-1.055297), (31710,-1.259618), (31711,-1.242375), (31712,-1.421149), (31713,-1.467076), (31714,-1.204116), (31715,-0.949980), (31716,-1.100884), (31717,-1.171431), (31718,-1.222004), (31719,-1.046833), (31720,-1.202846), (31721,-1.239020), (31722,-1.003000), (31723,-0.721924), (31724,-0.883975), (31725,-0.954987), (31726,-1.127722), (31727,-1.101189), (31728,-1.293433), (31729,-1.323568), (31730,-1.108915), (31731,-0.842703), (31732,-0.954589), (31733,-1.037676), (31734,-1.094288), (31735,-0.925620), (31736,-1.000812), (31737,-1.070428), (31738,-1.213900), (31739,-0.553332), (31740,-0.722816), (31741,-0.785931), (31742,-0.921971), (31743,-0.959074), (31744,-1.059348), (31745,-1.125249), (31746,-1.252464), (31747,-0.609546), (31748,-0.755341), (31749,-0.830068), (31750,-0.970288), (31751,-0.742629), (31752,-1.030559), (31753,-1.067662), (31754,-1.218566), (31755,-0.556140), (31756,-0.683819), (31757,-0.741824), (31758,-0.904340), (31759,-0.901032), (31760,-1.089096), (31761,-1.138740), (31762,-1.264097), (31763,-0.611425), (31764,-0.746536), (31765,-0.824979), (31766,-0.970309), (31767,-0.721283), (31768,-1.004568), (31769,-1.199134), (31770,-0.922703), (31771,-0.650452), (31772,-0.735398), (31773,-0.888625), (31774,-0.852802), (31775,-1.026931), (31776,-1.108625), (31777,-1.247916), (31778,-0.983562), (31779,-0.721530), (31780,-0.757704), (31781,-0.916505), (31782,-0.748765), (31783,-0.842536), (31784,-1.139756), (31785,-1.287408), (31786,-0.641240), (31787,-0.783318), (31788,-0.824601), (31789,-0.995479), (31790,-1.004712), (31791,-1.149577), (31792,-1.189932), (31793,-1.354771), (31794,-0.672371), (31795,-0.787973), (31796,-0.885925), (31797,-1.027539), (31798,-0.781300), (31799,-0.958680), (31800,-1.033871), (31801,-1.186169), (31802,-0.911131), (31803,-0.698336), (31804,-0.725220), (31805,-0.862653), (31806,-0.842159), (31807,-1.050196), (31808,-1.132819), (31809,-1.288368), (31810,-1.021227), (31811,-0.761982), (31812,-0.795833), (31813,-0.942557), (31814,-0.778998), (31815,-0.817030), (31816,-0.934490), (31817,-1.118373), (31818,-0.842871), (31819,-0.620785), (31820,-0.692725), (31821,-0.854313), (31822,-0.823599), (31823,-0.983329), (31824,-1.056662), (31825,-1.205708), (31826,-0.907446), (31827,-0.677000), (31828,-0.761481), (31829,-0.925855), (31830,-0.773909), (31831,-0.818443), (31832,-1.004649), (31833,-1.156018), (31834,-0.856826), (31835,-0.598511), (31836,-0.671379), (31837,-0.833895), (31838,-0.784138), (31839,-0.986136), (31840,-1.023704), (31841,-1.202477), (31842,-0.925117), (31843,-0.673769), (31844,-0.736418), (31845,-0.885000), (31846,-0.742344), (31847,-0.801277), (31848,-1.075272), (31849,-1.113304), (31850,-0.876355), (31851,-0.594815), (31852,-0.750828), (31853,-0.802330), (31854,-0.995503), (31855,-0.972222), (31856,-1.130558), (31857,-1.185776), (31858,-0.957187), (31859,-0.641739), (31860,-0.834912), (31861,-0.891058), (31862,-0.981114), (31863,-0.788756), (31864,-1.189558), (31865,-1.346965), (31866,-0.674784), (31867,-0.821508), (31868,-0.884623), (31869,-1.034598), (31870,-1.055908), (31871,-1.214244), (31872,-1.498457), (31873,-1.643787), (31874,-0.957208), (31875,-1.086280), (31876,-1.181445), (31877,-1.350000), (31878,-1.142314), (31879,-1.278354), (31880,-1.385595), (31881,-1.421769), (31882,-1.179246), (31883,-0.903744), (31884,-1.062544), (31885,-1.103363), (31886,-1.269131), (31887,-1.257926), (31888,-1.436236), (31889,-1.500744), (31890,-1.250788), (31891,-0.953920), (31892,-1.128977), (31893,-1.177692), (31894,-1.248239), (31895,-1.089789), (31896,-1.252770), (31897,-1.318207), (31898,-1.430558), (31899,-0.796001), (31900,-0.969666), (31901,-1.033709), (31902,-1.149312), (31903,-1.184557), (31904,-1.319203), (31905,-1.340513), (31906,-1.496526), (31907,-0.824811), (31908,-0.998474), (31909,-1.062518), (31910,-1.210171), (31911,-0.956964), (31912,-1.289950), (31913,-1.327053), (31914,-1.110542), (31915,-0.849903), (31916,-0.987801), (31917,-1.060671), (31918,-1.249198), (31919,-1.238923), (31920,-1.394936), (31921,-1.476166), (31922,-1.220637), (31923,-0.957676), (31924,-1.130411), (31925,-1.168908), (31926,-1.196720), (31927,-1.024801), (31928,-1.457653), (31929,-1.482679), (31930,-1.243407), (31931,-0.970227), (31932,-1.147143), (31933,-1.195394), (31934,-1.397857), (31935,-1.383400), (31936,-1.551955), (31937,-1.587200), (31938,-1.355825), (31939,-1.050595), (31940,-1.228905), (31941,-1.238138), (31942,-1.324941), (31943,-1.158131), (31944,-1.338762), (31945,-1.342422), (31946,-1.107795), (31947,-0.859698), (31948,-1.003170), (31949,-1.065820), (31950,-1.255742), (31951,-1.246859), (31952,-1.389403), (31953,-1.466452), (31954,-1.224393), (31955,-0.935421), (31956,-1.104905), (31957,-1.175916), (31958,-1.219057), (31959,-1.078723), (31960,-1.279792), (31961,-1.328971), (31962,-1.478947), (31963,-0.822094), (31964,-0.960922), (31965,-0.966438), (31966,-1.130349), (31967,-1.168845), (31968,-1.359231), (31969,-1.402837), (31970,-1.521690), (31971,-0.824427), (31972,-1.001807), (31973,-1.061206), (31974,-1.208858), (31975,-1.008140), (31976,-1.160437), (31977,-1.187785), (31978,-1.325683), (31979,-0.643285), (31980,-0.778860), (31981,-0.820607), (31982,-0.989627), (31983,-1.025336), (31984,-1.190175), (31985,-1.240748), (31986,-1.406051), (31987,-0.712504), (31988,-0.916361), (31989,-0.955786), (31990,-1.121554), (31991,-0.897146), (31992,-1.115866), (31993,-1.174336), (31994,-1.327098), (31995,-0.646091), (31996,-0.784454), (31997,-0.852214), (31998,-0.961777), (31999,-1.011886), (32000,-1.092187), (32001,-1.130218), (32002,-1.283909), (32003,-0.646566), (32004,-0.758917), (32005,-0.836431), (32006,-0.991051), (32007,-0.745276), (32008,-1.073618), (32009,-1.098179), (32010,-1.254192), (32011,-0.564361), (32012,-0.723626), (32013,-0.829938), (32014,-0.978984), (32015,-0.977534), (32016,-1.154914), (32017,-1.188765), (32018,-1.353139), (32019,-0.693965), (32020,-0.871810), (32021,-0.911699), (32022,-1.031947), (32023,-0.807539), (32024,-1.103830), (32025,-1.249624), (32026,-0.930924), (32027,-0.706052), (32028,-0.762199), (32029,-0.908923), (32030,-0.894002), (32031,-1.027719), (32032,-1.112201), (32033,-1.296549), (32034,-1.018724), (32035,-0.772949), (32036,-0.818413), (32037,-0.965601), (32038,-0.825731), (32039,-0.925076), (32040,-1.103386), (32041,-1.248715), (32042,-0.967175), (32043,-0.714433), (32044,-0.772903), (32045,-0.927523), (32046,-0.940472), (32047,-1.079763), (32048,-1.118259), (32049,-1.279382), (32050,-1.023853), (32051,-0.801304), (32052,-0.843052), (32053,-0.975840), (32054,-0.825752), (32055,-0.904194), (32056,-1.031874), (32057,-1.246878), (32058,-0.964873), (32059,-0.680545), (32060,-0.724616), (32061,-0.907105), (32062,-0.908907), (32063,-1.084893), (32064,-1.124318), (32065,-1.277080), (32066,-1.002507), (32067,-0.806433), (32068,-0.870012), (32069,-1.019058), (32070,-0.836920), (32071,-0.907466), (32072,-1.030965), (32073,-1.222745), (32074,-0.975112), (32075,-0.701932), (32076,-0.766440), (32077,-0.948465), (32078,-0.943764), (32079,-1.122537), (32080,-1.169859), (32081,-1.315653), (32082,-1.035506), (32083,-0.791590), (32084,-0.822190), (32085,-0.974952), (32086,-0.829508), (32087,-0.918170), (32088,-1.037488), (32089,-1.162381), (32090,-0.907316), (32091,-0.698237), (32092,-0.759029), (32093,-0.910397), (32094,-0.907089), (32095,-1.069141), (32096,-1.143403), (32097,-1.283159), (32098,-1.027630), (32099,-0.746090), (32100,-0.814778), (32101,-0.996339), (32102,-0.855075), (32103,-0.933054), (32104,-1.181966), (32105,-1.316148), (32106,-0.606344), (32107,-0.760499), (32108,-0.825936), (32109,-0.992168), (32110,-0.996756), (32111,-1.144409), (32112,-1.217278), (32113,-1.342635), (32114,-0.694144), (32115,-0.839009), (32116,-0.895156), (32117,-1.034912), (32118,-0.799356), (32119,-0.951654), (32120,-1.287891), (32121,-1.432757), (32122,-0.769402), (32123,-0.929131), (32124,-0.992245), (32125,-1.164516), (32126,-1.170033), (32127,-1.310718), (32128,-1.344570), (32129,-1.495009), (32130,-1.233442), (32131,-0.965836), (32132,-0.977392), (32133,-1.157094), (32134,-1.012115), (32135,-1.080339), (32136,-1.231708), (32137,-1.316653), (32138,-1.448513), (32139,-0.798164), (32140,-0.941636), (32141,-1.012182), (32142,-1.180273), (32143,-1.200189), (32144,-1.345519), (32145,-1.386338), (32146,-1.546067), (32147,-0.872029), (32148,-0.998779), (32149,-1.068396), (32150,-1.224874), (32151,-0.996286), (32152,-1.275855), (32153,-1.352904), (32154,-1.494983), (32155,-0.797255), (32156,-0.963023), (32157,-1.004306), (32158,-1.119909), (32159,-1.147257), (32160,-1.325102), (32161,-1.404473), (32162,-1.582782), (32163,-0.867869), (32164,-1.010412), (32165,-1.067023), (32166,-1.210031), (32167,-0.974940), (32168,-1.374813), (32169,-1.423992), (32170,-1.173108), (32171,-0.893890), (32172,-1.058729), (32173,-1.118592), (32174,-1.295043), (32175,-1.288484), (32176,-1.433349), (32177,-1.503895), (32178,-1.249760), (32179,-0.961717), (32180,-1.118195), (32181,-1.200353), (32182,-1.268113), (32183,-1.120347), (32184,-1.315378), (32185,-1.347371), (32186,-1.519177), (32187,-0.825165), (32188,-0.971424), (32189,-1.032681), (32190,-1.178011), (32191,-1.206288), (32192,-1.346509), (32193,-1.391973), (32194,-1.534980), (32195,-0.884166), (32196,-1.009523), (32197,-1.088895), (32198,-1.250947), (32199,-1.047906), (32200,-1.219247), (32201,-1.297690), (32202,-1.449988), (32203,-0.757834), (32204,-0.908738), (32205,-0.966743), (32206,-1.135298), (32207,-1.157537), (32208,-1.295899), (32209,-1.341363), (32210,-1.492267), (32211,-0.821480), (32212,-0.977029), (32213,-1.052220), (32214,-1.206840), (32215,-0.948060), (32216,-1.287084), (32217,-1.339515), (32218,-1.474626), (32219,-0.821955), (32220,-0.969142), (32221,-1.035508), (32222,-1.196167), (32223,-1.225373), (32224,-1.375813), (32225,-1.439391), (32226,-1.565213), (32227,-0.878169), (32228,-1.007706), (32229,-1.078717), (32230,-1.222189), (32231,-0.998245), (32232,-1.130105), (32233,-1.210406), (32234,-1.381748), (32235,-0.688200), (32236,-0.841427), (32237,-0.896645), (32238,-1.019215), (32239,-1.043312), (32240,-1.186784), (32241,-1.242931), (32242,-1.428672), (32243,-0.748130), (32244,-0.895783), (32245,-0.977013), (32246,-1.126987), (32247,-0.881213), (32248,-1.197477), (32249,-1.255018), (32250,-1.377123), (32251,-0.735599), (32252,-0.864672), (32253,-0.903633), (32254,-1.074510), (32255,-1.080027), (32256,-1.212351), (32257,-1.294974), (32258,-1.431943), (32259,-0.750473), (32260,-0.900448), (32261,-0.977962), (32262,-1.109821), (32263,-0.884020), (32264,-1.119927), (32265,-1.194189), (32266,-1.401297), (32267,-0.720756), (32268,-0.891168), (32269,-0.946851), (32270,-1.097290), (32271,-1.099091), (32272,-1.246744), (32273,-1.303820), (32274,-1.426854), (32275,-0.787188), (32276,-0.939950), (32277,-0.999813), (32278,-1.145608), (32279,-0.906801), (32280,-1.048415), (32281,-1.193745), (32282,-0.912669), (32283,-1.077508), (32284,-0.765775), (32285,-0.891132), (32286,-0.906403), (32287,-1.073100), (32288,-1.158046), (32289,-1.296873), (32290,-1.030661), (32291,-1.203860), (32292,-0.859613), (32293,-1.002156), (32294,-0.851603), (32295,-1.017371), (32296,-1.117645), (32297,-1.269478), (32298,-1.046928), (32299,-0.777464), (32300,-0.845224), (32301,-0.991483), (32302,-0.965879), (32303,-1.151155), (32304,-1.170607), (32305,-1.340091), (32306,-1.056693), (32307,-0.814170), (32308,-0.911192), (32309,-1.020756), (32310,-0.874384), (32311,-0.901268), (32312,-1.183159), (32313,-1.370758), (32314,-1.071567), (32315,-0.831831), (32316,-0.876830), (32317,-1.003580), (32318,-1.023497), (32319,-1.189729), (32320,-1.233799), (32321,-1.402818), (32322,-1.118955), (32323,-0.873181), (32324,-0.923289), (32325,-1.076051), (32326,-0.916673), (32327,-1.000225), (32328,-1.126046), (32329,-1.284847), (32330,-1.004700), (32331,-0.756603), (32332,-0.778377), (32333,-0.928352), (32334,-0.955701), (32335,-1.129829), (32336,-1.198053), (32337,-1.339667), (32338,-1.069739), (32339,-0.819320), (32340,-0.874538), (32341,-1.048202), (32342,-0.899507), (32343,-0.971911), (32344,-1.031310), (32345,-1.183143), (32346,-0.903925), (32347,-1.027423), (32348,-0.697575), (32349,-0.848015), (32350,-0.839597), (32351,-1.017906), (32352,-1.093562), (32353,-1.232854), (32354,-0.954100), (32355,-1.122655), (32356,-0.769582), (32357,-0.921415), (32358,-0.782010), (32359,-0.942204), (32360,-1.238030), (32361,-1.277455), (32362,-1.053512), (32363,-0.768720), (32364,-0.901044), (32365,-0.953940), (32366,-1.150364), (32367,-1.107574), (32368,-1.291922), (32369,-1.333669), (32370,-1.155247), (32371,-0.818431), (32372,-0.967942), (32373,-1.062642), (32374,-1.142943), (32375,-0.985887), (32376,-1.140971), (32377,-1.313706), (32378,-1.007547), (32379,-0.770598), (32380,-0.833713), (32381,-1.000410), (32382,-0.987812), (32383,-1.172624), (32384,-1.513970), (32385,-1.542248), (32386,-1.287648), (32387,-1.007965), (32388,-1.145863), (32389,-1.192256), (32390,-1.286492), (32391,-1.129900), (32392,-1.360233), (32393,-1.388046), (32394,-1.137162), (32395,-0.856550), (32396,-0.997235), (32397,-1.098903), (32398,-1.284644), (32399,-1.266472), (32400,-1.422021), (32401,-1.482813), (32402,-1.226355), (32403,-0.927164), (32404,-1.080390), (32405,-1.122138), (32406,-1.205225), (32407,-1.065356), (32408,-1.095956), (32409,-1.252898), (32410,-1.311832), (32411,-1.040510), (32412,-0.774298), (32413,-0.911267), (32414,-0.972059), (32415,-1.165232), (32416,-1.154492), (32417,-1.283100), (32418,-1.358292), (32419,-1.097653), (32420,-0.825867), (32421,-0.972591), (32422,-1.040350), (32423,-1.128547), (32424,-1.149857), (32425,-1.280788), (32426,-0.937470), (32427,-1.101844), (32428,-0.834703), (32429,-0.950305), (32430,-1.058940), (32431,-1.248397), (32432,-1.191672), (32433,-1.317029), (32434,-1.011799), (32435,-1.160845), (32436,-0.925754), (32437,-1.063187), (32438,-1.015288), (32439,-1.168514), (32440,-1.305483), (32441,-1.483328), (32442,-1.138616), (32443,-1.299274), (32444,-0.998225), (32445,-1.161206), (32446,-1.232217), (32447,-1.410526), (32448,-1.388638), (32449,-1.568341), (32450,-1.217126), (32451,-1.351772), (32452,-1.069303), (32453,-1.193731), (32454,-1.113316), (32455,-1.268865), (32456,-1.188915), (32457,-1.375121), (32458,-1.032267), (32459,-1.186423), (32460,-0.937397), (32461,-1.052999), (32462,-1.137016), (32463,-1.297210), (32464,-1.294366), (32465,-1.417400), (32466,-1.127034), (32467,-1.303950), (32468,-1.034486), (32469,-1.174242), (32470,-1.169540), (32471,-1.303258), (32472,-1.145738), (32473,-1.318008), (32474,-1.374155), (32475,-1.122807), (32476,-0.851485), (32477,-1.001460), (32478,-1.059930), (32479,-1.202008), (32480,-1.195449), (32481,-1.376545), (32482,-1.430834), (32483,-1.168338), (32484,-0.866359), (32485,-1.046527), (32486,-1.067836), (32487,-1.124448), (32488,-0.971573), (32489,-1.152204), (32490,-1.232040), (32491,-0.956538), (32492,-0.708441), (32493,-0.867706), (32494,-0.912705), (32495,-1.096124), (32496,-1.082132), (32497,-1.252545), (32498,-1.279429), (32499,-1.043873), (32500,-0.797170), (32501,-0.927172), (32502,-0.971242), (32503,-1.027389), (32504,-0.917711), (32505,-1.094627), (32506,-1.087138), (32507,-0.872485), (32508,-0.605344), (32509,-0.740920), (32510,-0.798460), (32511,-0.949828), (32512,-1.015265), (32513,-1.173601), (32514,-1.202343), (32515,-0.965394), (32516,-0.688034), (32517,-0.825003), (32518,-0.909020), (32519,-0.967489), (32520,-0.980438), (32521,-1.135523), (32522,-1.188883), (32523,-0.984449), (32524,-0.706624), (32525,-0.868676), (32526,-0.920178), (32527,-1.081765), (32528,-1.104469), (32529,-1.251657), (32530,-1.307804), (32531,-1.045772), (32532,-0.761444), (32533,-0.919780), (32534,-0.969889), (32535,-1.035326), (32536,-1.131419), (32537,-1.163413), (32538,-1.302704), (32539,-0.637491), (32540,-0.773067), (32541,-0.872877), (32542,-1.001949), (32543,-1.007466), (32544,-1.173234), (32545,-1.213124), (32546,-1.360776), (32547,-0.665836), (32548,-0.802340), (32549,-0.910046), (32550,-1.062344), (32551,-0.809602), (32552,-1.082668), (32553,-1.142531), (32554,-1.325485), (32555,-0.658878), (32556,-0.763333), (32557,-0.834808), (32558,-1.014975), (32559,-0.999590), (32560,-1.160713), (32561,-1.231724), (32562,-1.360797), (32563,-0.697442), (32564,-0.849739), (32565,-0.868726), (32566,-1.035423), (32567,-0.824486), (32568,-1.071076), (32569,-1.126758), (32570,-1.263727), (32571,-0.578541), (32572,-0.735948), (32573,-0.795347), (32574,-0.934174), (32575,-0.949910), (32576,-1.104065), (32577,-1.178792), (32578,-1.348740), (32579,-0.643581), (32580,-0.802845), (32581,-0.899403), (32582,-1.039624), (32583,-0.794314), (32584,-1.053445), (32585,-1.076613), (32586,-1.222872), (32587,-0.567878), (32588,-0.704383), (32589,-0.762852), (32590,-0.912363), (32591,-0.935066), (32592,-1.103156), (32593,-1.163019), (32594,-1.313459), (32595,-0.650104), (32596,-0.803795), (32597,-0.848329), (32598,-1.006665), (32599,-0.775755), (32600,-1.021415), (32601,-1.069202), (32602,-1.224750), (32603,-0.552106), (32604,-0.710906), (32605,-0.765659), (32606,-0.936537), (32607,-0.942518), (32608,-1.080416), (32609,-1.159788), (32610,-1.331130), (32611,-0.648266), (32612,-0.785235), (32613,-0.847885), (32614,-1.030839), (32615,-0.759982), (32616,-1.139882), (32617,-1.205319), (32618,-0.979518), (32619,-0.686365), (32620,-0.785710), (32621,-0.848824), (32622,-1.005302), (32623,-0.971802), (32624,-1.101803), (32625,-1.173743), (32626,-0.971167), (32627,-0.701703), (32628,-0.849356), (32629,-0.918044), (32630,-0.983017), (32631,-0.835715), (32632,-1.261135), (32633,-1.333075), (32634,-1.057573), (32635,-0.771388), (32636,-0.925078), (32637,-0.999805), (32638,-1.177650), (32639,-1.145543), (32640,-1.124119), (32641,-0.803097), (32642,-0.923344), (32643,-0.642268), (32644,-0.813610), (32645,-0.772678), (32646,-0.910576), (32647,-0.760952), (32648,-0.917429), (32649,-0.722285), (32650,-0.746382), (32651,-0.918653), (32652,-0.642222), (32653,-0.797306), (32654,-0.852988), (32655,-1.002034), (32656,-0.978288), (32657,-0.732514), (32658,-0.796557), (32659,-0.947926), (32660,-0.668243), (32661,-0.748080), (32662,-0.825593), (32663,-0.999722), (32664,-0.799933), (32665,-0.953624), (32666,-0.614950), (32667,-0.755171), (32668,-0.502429), (32669,-0.663552), (32670,-0.704371), (32671,-0.865493), (32672,-0.861256), (32673,-1.014482), (32674,-0.688351), (32675,-0.833216), (32676,-0.563288), (32677,-0.717908), (32678,-0.702523), (32679,-0.865039), (32680,-0.872879), (32681,-0.595519), (32682,-0.674890), (32683,-0.807679), (32684,-0.563298), (32685,-0.738356), (32686,-0.805651), (32687,-0.977921), (32688,-0.970897), (32689,-0.728839), (32690,-0.774302), (32691,-0.916381), (32692,-0.626944), (32693,-0.701206), (32694,-0.745276), (32695,-0.888748), (32696,-1.004815), (32697,-0.769724), (32698,-0.840735), (32699,-0.997678), (32700,-0.707776), (32701,-0.902343), (32702,-0.943161), (32703,-1.090349), (32704,-1.067532), (32705,-0.828261), (32706,-0.853751), (32707,-1.019983), (32708,-0.732404), (32709,-0.803415), (32710,-0.844234), (32711,-1.017434), (32712,-0.915188), (32713,-0.706573), (32714,-0.741354), (32715,-0.886684), (32716,-0.605143), (32717,-0.747222), (32718,-0.797330), (32719,-0.928261), (32720,-0.920772), (32721,-0.715873), (32722,-0.759944), (32723,-0.902487), (32724,-0.633952), (32725,-0.700782), (32726,-0.738814), (32727,-0.917588), (32728,-0.789795), (32729,-0.922584), (32730,-0.603419), (32731,-0.760361), (32732,-0.476498), (32733,-0.660846), (32734,-0.732321), (32735,-0.860465), (32736,-0.825107), (32737,-0.990410), (32738,-0.656846), (32739,-0.828652), (32740,-0.552686), (32741,-0.713808), (32742,-0.685882), (32743,-0.838179), (32744,-0.705277), (32745,-0.866864), (32746,-0.519830), (32747,-0.675844), (32748,-0.372936), (32749,-0.533130), (32750,-0.606464), (32751,-0.754581), (32752,-0.751272), (32753,-0.897531), (32754,-0.547710), (32755,-0.726019), (32756,-0.453304), (32757,-0.599099), (32758,-0.558631), (32759,-0.690026), (32760,-0.617043), (32761,-0.750761), (32762,-0.399546), (32763,-0.543018), (32764,-0.253582), (32765,-0.423530), (32766,-0.495470), (32767,-0.647767), (32768,-0.652355), (32769,-0.821374), (32770,-0.474340), (32771,-0.632676), (32772,-0.316763), (32773,-0.485318), (32774,-0.457391), (32775,-0.643597), (32776,-0.617064), (32777,-0.782367), (32778,-0.411644), (32779,-0.559296), (32780,-0.300516), (32781,-0.459781), (32782,-0.534507), (32783,-0.694701), (32784,-0.658414), (32785,-0.821859), (32786,-0.487831), (32787,-0.651741), (32788,-0.374381), (32789,-0.525749), (32790,-0.519654), (32791,-0.638972), (32792,-0.821462), (32793,-0.865067), (32794,-0.587707), (32795,-0.358190), (32796,-0.532783), (32797,-0.598685), (32798,-0.770955), (32799,-0.723985), (32800,-0.879069), (32801,-0.951938), (32802,-0.689906), (32803,-0.393966), (32804,-0.537438), (32805,-0.612165), (32806,-0.695718), (32807,-0.540055), (32808,-0.745769), (32809,-0.802381), (32810,-0.580760), (32811,-0.281569), (32812,-0.418538), (32813,-0.442635), (32814,-0.631627), (32815,-0.626461), (32816,-0.796409), (32817,-0.852556), (32818,-0.587738), (32819,-0.318274), (32820,-0.487758), (32821,-0.533686), (32822,-0.585653), (32823,-0.451357), (32824,-0.729068), (32825,-0.810298), (32826,-0.564523), (32827,-0.269977), (32828,-0.423203), (32829,-0.460306), (32830,-0.667878), (32831,-0.621372), (32832,-0.784353), (32833,-0.835390), (32834,-0.595654), (32835,-0.326191), (32836,-0.486385), (32837,-0.516056), (32838,-0.602395), (32839,-0.444874), (32840,-0.728624), (32841,-0.748076), (32842,-0.555718), (32843,-0.248166), (32844,-0.389315), (32845,-0.457075), (32846,-0.639100), (32847,-0.608851), (32848,-0.775548), (32849,-0.842843), (32850,-0.602642), (32851,-0.306238), (32852,-0.458071), (32853,-0.481703), (32854,-0.577332), (32855,-0.426779), (32856,-0.749546), (32857,-0.820093), (32858,-0.600330), (32859,-0.302067), (32860,-0.465513), (32861,-0.503545), (32862,-0.704149), (32863,-0.653463), (32864,-0.819230), (32865,-0.876771), (32866,-0.631461), (32867,-0.379184), (32868,-0.521727), (32869,-0.553720), (32870,-0.646562), (32871,-0.503441), (32872,-0.758856), (32873,-0.428544), (32874,-0.565978), (32875,-0.322061), (32876,-0.451134), (32877,-0.523074), (32878,-0.685125), (32879,-0.673921), (32880,-0.830399), (32881,-0.521917), (32882,-0.663067), (32883,-0.369914), (32884,-0.546830), (32885,-0.530516), (32886,-0.666091), (32887,-0.537834), (32888,-0.973009), (32889,-0.608324), (32890,-0.757370), (32891,-0.461430), (32892,-0.610940), (32893,-0.673126), (32894,-0.823565), (32895,-0.849520), (32896,-0.855037), (32897,-0.892140), (32898,-0.679809), (32899,-0.534830), (32900,-0.687127), (32901,-0.723766), (32902,-0.786416), (32903,-0.505804), (32904,-0.756574), (32905,-0.802967), (32906,-0.592494), (32907,-0.611482), (32908,-0.756812), (32909,-0.806456), (32910,-0.979191), (32911,-0.679535), (32912,-0.823936), (32913,-0.858252), (32914,-0.653818), (32915,-0.460531), (32916,-0.620260), (32917,-0.676872), (32918,-0.768785), (32919,-0.454730), (32920,-0.699926), (32921,-0.722165), (32922,-0.486145), (32923,-0.493520), (32924,-0.676010), (32925,-0.763278), (32926,-0.915111), (32927,-0.629390), (32928,-0.798874), (32929,-0.847125), (32930,-0.625968), (32931,-0.444294), (32932,-0.622603), (32933,-0.678750), (32934,-0.761374), (32935,-0.451034), (32936,-0.795633), (32937,-0.577263), (32938,-0.631552), (32939,-0.782921), (32940,-0.788438), (32941,-0.965354), (32942,-1.008495), (32943,-1.139890), (32944,-0.879716), (32945,-0.628832), (32946,-0.691947), (32947,-0.873507), (32948,-0.705768), (32949,-0.796752), (32950,-0.865905), (32951,-1.029815), (32952,-0.784505), (32953,-0.943770), (32954,-0.602309), (32955,-0.727202), (32956,-0.732254), (32957,-0.877120), (32958,-0.982503), (32959,-1.124117), (32960,-0.827249), (32961,-0.991623), (32962,-0.621364), (32963,-0.794564), (32964,-0.608244), (32965,-0.782373), (32966,-0.754447), (32967,-0.884448), (32968,-0.698594), (32969,-0.856465), (32970,-0.481561), (32971,-0.651974), (32972,-0.650988), (32973,-0.754049), (32974,-0.855717), (32975,-0.996402), (32976,-0.726009), (32977,-0.882022), (32978,-0.556355), (32979,-0.706330), (32980,-0.582253), (32981,-0.695533), (32982,-0.631376), (32983,-0.802718), (32984,-0.682821), (32985,-0.812358), (32986,-0.482975), (32987,-0.650136), (32988,-0.664943), (32989,-0.786120), (32990,-0.871530), (32991,-1.022898), (32992,-0.705592), (32993,-0.860211), (32994,-0.561949), (32995,-0.705421), (32996,-0.567874), (32997,-0.696947), (32998,-0.705715), (32999,-0.821318), (33000,-0.541171), (33001,-0.703222), (33002,-0.397528), (33003,-0.514524), (33004,-0.505642), (33005,-0.654688), (33006,-0.786083), (33007,-0.924910), (33008,-0.643370), (33009,-0.739928), (33010,-0.390106), (33011,-0.563771), (33012,-0.412289), (33013,-0.579914), (33014,-0.568245), (33015,-0.698247), (33016,-0.567203), (33017,-0.695346), (33018,-0.344132), (33019,-0.507577), (33020,-0.528422), (33021,-0.667250), (33022,-0.728970), (33023,-0.892880), (33024,-0.646641), (33025,-0.823092), (33026,-0.469091), (33027,-0.591661), (33028,-0.450397), (33029,-0.606411), (33030,-0.558976), (33031,-0.723814), (33032,-0.621104), (33033,-0.787337), (33034,-0.462598), (33035,-0.604212), (33036,-0.612981), (33037,-0.731370), (33038,-0.843721), (33039,-1.002521), (33040,-0.734916), (33041,-0.884891), (33042,-0.554114), (33043,-0.670181), (33044,-0.504299), (33045,-0.667744), (33046,-0.613342), (33047,-0.787006), (33048,-0.725636), (33049,-0.790608), (33050,-0.530435), (33051,-0.532236), (33052,-0.697075), (33053,-0.756938), (33054,-0.944537), (33055,-0.646274), (33056,-0.814364), (33057,-0.855183), (33058,-0.643317), (33059,-0.506234), (33060,-0.614405), (33061,-0.686344), (33062,-0.729486), (33063,-0.441907), (33064,-0.610461), (33065,-0.677292), (33066,-0.440343), (33067,-0.430532), (33068,-0.585152), (33069,-0.591133), (33070,-0.792203), (33071,-0.561757), (33072,-0.702906), (33073,-0.784136), (33074,-0.538826), (33075,-0.355294), (33076,-0.526171), (33077,-0.546087), (33078,-0.614776), (33079,-0.347635), (33080,-0.716387), (33081,-0.761386), (33082,-0.491458), (33083,-0.510445), (33084,-0.711514), (33085,-0.739327), (33086,-0.899521), (33087,-0.595685), (33088,-0.786535), (33089,-0.801342), (33090,-0.598301), (33091,-0.436136), (33092,-0.596330), (33093,-0.641794), (33094,-0.719307), (33095,-0.453560), (33096,-0.750315), (33097,-0.762800), (33098,-0.541643), (33099,-0.537406), (33100,-0.695277), (33101,-0.754676), (33102,-0.942275), (33103,-0.648658), (33104,-0.814890), (33105,-0.843167), (33106,-0.622011), (33107,-0.464955), (33108,-0.621433), (33109,-0.715668), (33110,-0.739765), (33111,-0.478663), (33112,-0.719214), (33113,-0.760497), (33114,-0.505897), (33115,-0.508628), (33116,-0.662783), (33117,-0.675732), (33118,-0.878659), (33119,-0.633350), (33120,-0.782860), (33121,-0.823679), (33122,-0.568150), (33123,-0.423171), (33124,-0.614950), (33125,-0.644157), (33126,-0.700304), (33127,-0.440594), (33128,-0.802843), (33129,-0.465099), (33130,-0.625293), (33131,-0.594115), (33132,-0.738051), (33133,-0.842970), (33134,-1.011990), (33135,-0.701186), (33136,-0.859057), (33137,-0.523171), (33138,-0.665250), (33139,-0.519806), (33140,-0.666065), (33141,-0.633494), (33142,-0.778824), (33143,-0.537694), (33144,-0.706713), (33145,-0.731275), (33146,-0.510583), (33147,-0.494269), (33148,-0.642850), (33149,-0.717113), (33150,-0.866159), (33151,-0.581367), (33152,-0.780114), (33153,-0.911509), (33154,-0.566332), (33155,-0.700515), (33156,-0.572257), (33157,-0.702259), (33158,-0.672939), (33159,-0.820127), (33160,-0.670503), (33161,-0.836271), (33162,-0.499920), (33163,-0.621096), (33164,-0.621504), (33165,-0.803065), (33166,-0.879649), (33167,-1.012438), (33168,-0.739258), (33169,-0.885517), (33170,-0.529193), (33171,-0.685671), (33172,-0.552304), (33173,-0.715750), (33174,-0.671101), (33175,-0.815038), (33176,-0.679813), (33177,-0.821892), (33178,-0.490650), (33179,-0.588602), (33180,-0.646607), (33181,-0.745952), (33182,-0.840652), (33183,-0.983195), (33184,-0.736027), (33185,-0.895292), (33186,-0.525033), (33187,-0.693588), (33188,-0.579265), (33189,-0.699513), (33190,-0.643717), (33191,-0.797407), (33192,-0.782022), (33193,-0.526029), (33194,-0.582176), (33195,-0.721932), (33196,-0.756712), (33197,-0.913655), (33198,-0.932642), (33199,-1.106771), (33200,-0.831269), (33201,-0.589210), (33202,-0.659757), (33203,-0.807874), (33204,-0.658250), (33205,-0.756201), (33206,-0.771937), (33207,-0.953033), (33208,-0.714691), (33209,-0.865595), (33210,-0.522277), (33211,-0.678290), (33212,-0.696813), (33213,-0.837498), (33214,-0.915941), (33215,-1.088676), (33216,-0.807135), (33217,-0.950607), (33218,-0.611470), (33219,-0.765625), (33220,-0.610427), (33221,-0.750648), (33222,-0.739907), (33223,-0.893598), (33224,-0.587440), (33225,-0.749027), (33226,-0.435901), (33227,-0.584018), (33228,-0.582568), (33229,-0.709782), (33230,-0.785438), (33231,-0.938200), (33232,-0.666878), (33233,-0.796880), (33234,-0.474928), (33235,-0.609111), (33236,-0.444623), (33237,-0.602494), (33238,-0.584322), (33239,-0.737084), (33240,-0.704048), (33241,-0.879106), (33242,-0.569231), (33243,-0.674150), (33244,-0.690351), (33245,-0.807346), (33246,-0.883467), (33247,-1.057595), (33248,-0.764442), (33249,-0.909308), (33250,-0.608723), (33251,-0.748944), (33252,-0.584920), (33253,-0.752082), (33254,-0.756670), (33255,-0.883885), (33256,-0.925168), (33257,-0.640840), (33258,-0.376486), (33259,-0.449355), (33260,-0.631380), (33261,-0.601596), (33262,-0.768757), (33263,-0.839303), (33264,-1.002748), (33265,-0.712847), (33266,-0.461499), (33267,-0.493492), (33268,-0.649505), (33269,-0.517997), (33270,-0.575537), (33271,-0.608460), (33272,-0.562882), (33273,-0.726328), (33274,-0.412737), (33275,-0.562247), (33276,-0.545004), (33277,-0.705663), (33278,-0.778067), (33279,-0.951731), (33280,-0.630709), (33281,-0.788580), (33282,-0.434114), (33283,-0.604991), (33284,-0.465121), (33285,-0.617419), (33286,-0.604821), (33287,-0.706953), (33288,-0.904771), (33289,-0.655745), (33290,-0.401609), (33291,-0.451718), (33292,-0.596583), (33293,-0.562154), (33294,-0.780874), (33295,-0.851885), (33296,-1.017653), (33297,-0.715675), (33298,-0.439244), (33299,-0.480062), (33300,-0.642579), (33301,-0.515250), (33302,-0.610879), (33303,-0.641015), (33304,-0.551310), (33305,-0.593987), (33306,-0.757897), (33307,-0.352801), (33308,-0.507421), (33309,-0.560781), (33310,-0.714472), (33311,-0.462659), (33312,-0.629356), (33313,-0.730559), (33314,-0.912119), (33315,-0.343521), (33316,-0.466091), (33317,-0.528741), (33318,-0.645272), (33319,-0.338649), (33320,-0.580129), (33321,-0.716634), (33322,-0.361239), (33323,-0.505175), (33324,-0.541814), (33325,-0.678318), (33326,-0.743755), (33327,-0.845887), (33328,-0.581069), (33329,-0.759378), (33330,-0.423956), (33331,-0.584150), (33332,-0.440100), (33333,-0.610512), (33334,-0.569115), (33335,-0.679144), (33336,-0.694880), (33337,-0.758923), (33338,-0.521045), (33339,-0.538175), (33340,-0.714161), (33341,-0.746155), (33342,-0.907278), (33343,-0.603906), (33344,-0.777570), (33345,-0.848581), (33346,-0.634857), (33347,-0.424848), (33348,-0.572501), (33349,-0.620751), (33350,-0.688046), (33351,-0.447846), (33352,-0.581563), (33353,-0.731074), (33354,-0.384969), (33355,-0.533086), (33356,-0.532564), (33357,-0.679288), (33358,-0.746583), (33359,-0.903061), (33360,-0.624307), (33361,-0.766386), (33362,-0.441183), (33363,-0.599983), (33364,-0.474513), (33365,-0.574787), (33366,-0.574730), (33367,-0.755362), (33368,-0.540244), (33369,-0.613113), (33370,-0.784454), (33371,-0.365888), (33372,-0.522830), (33373,-0.588267), (33374,-0.728023), (33375,-0.431619), (33376,-0.603890), (33377,-0.673972), (33378,-0.806760), (33379,-0.268819), (33380,-0.422974), (33381,-0.471225), (33382,-0.597975), (33383,-0.232361), (33384,-0.647098), (33385,-0.420368), (33386,-0.446323), (33387,-0.601871), (33388,-0.592060), (33389,-0.762473), (33390,-0.796789), (33391,-0.947693), (33392,-0.664759), (33393,-0.438958), (33394,-0.490460), (33395,-0.645080), (33396,-0.487559), (33397,-0.588762), (33398,-0.611001), (33399,-0.790239), (33400,-0.533781), (33401,-0.664248), (33402,-0.346476), (33403,-0.516425), (33404,-0.517762), (33405,-0.640331), (33406,-0.736889), (33407,-0.866891), (33408,-0.715874), (33409,-0.865384), (33410,-0.529033), (33411,-0.679473), (33412,-0.561434), (33413,-0.716054), (33414,-0.687198), (33415,-0.815806), (33416,-0.642494), (33417,-0.798043), (33418,-0.470517), (33419,-0.603306), (33420,-0.618113), (33421,-0.761120), (33422,-0.854891), (33423,-1.008117), (33424,-0.747944), (33425,-0.865869), (33426,-0.542988), (33427,-0.694356), (33428,-0.553558), (33429,-0.705855), (33430,-0.686290), (33431,-0.860883), (33432,-0.727052), (33433,-0.875169), (33434,-0.548108), (33435,-0.719914), (33436,-0.673407), (33437,-0.822454), (33438,-0.908793), (33439,-1.044833), (33440,-0.796272), (33441,-0.946247), (33442,-0.606180), (33443,-0.724569), (33444,-0.564261), (33445,-0.718417), (33446,-0.706748), (33447,-0.869264), (33448,-0.972325), (33449,-0.666631), (33450,-0.412031), (33451,-0.483971), (33452,-0.651132), (33453,-0.648753), (33454,-0.818701), (33455,-0.881351), (33456,-1.037365), (33457,-0.767436), (33458,-0.503547), (33459,-0.552262), (33460,-0.672974), (33461,-0.535891), (33462,-0.599006), (33463,-0.678842), (33464,-1.019724), (33465,-0.725642), (33466,-0.475687), (33467,-0.545769), (33468,-0.725007), (33469,-0.714732), (33470,-0.880034), (33471,-0.928750), (33472,-1.106595), (33473,-0.821338), (33474,-0.612723), (33475,-0.634033), (33476,-0.774718), (33477,-0.606514), (33478,-0.685421), (33479,-0.719738), (33480,-0.903156), (33481,-0.629048), (33482,-0.398601), (33483,-0.466360), (33484,-0.633058), (33485,-0.594448), (33486,-0.790408), (33487,-0.835871), (33488,-0.961692), (33489,-0.693622), (33490,-0.476647), (33491,-0.529542), (33492,-0.691130), (33493,-0.543828), (33494,-0.620877), (33495,-0.657980), (33496,-1.094548), (33497,-0.819511), (33498,-0.566304), (33499,-0.613626), (33500,-0.789612), (33501,-0.737532), (33502,-0.916306), (33503,-0.971059), (33504,-1.149368), (33505,-0.903129), (33506,-0.649459), (33507,-0.685633), (33508,-0.838859), (33509,-0.681339), (33510,-0.765820), (33511,-0.829864), (33512,-0.972871), (33513,-0.657886), (33514,-0.444627), (33515,-0.560229), (33516,-0.716243), (33517,-0.670201), (33518,-0.849439), (33519,-0.903263), (33520,-1.041626), (33521,-0.756370), (33522,-0.512453), (33523,-0.548627), (33524,-0.726936), (33525,-0.580099), (33526,-0.624169), (33527,-0.677994), (33528,-0.747147), (33529,-0.510198), (33530,-0.661102), (33531,-0.316854), (33532,-0.464042), (33533,-0.495571), (33534,-0.619070), (33535,-0.677539), (33536,-0.755982), (33537,-0.492557), (33538,-0.670866), (33539,-0.313613), (33540,-0.480774), (33541,-0.321861), (33542,-0.519678), (33543,-0.457844), (33544,-0.776430), (33545,-0.481419), (33546,-0.661586), (33547,-0.300153), (33548,-0.455702), (33549,-0.481192), (33550,-0.620484), (33551,-0.715184), (33552,-0.855404), (33553,-0.587334), (33554,-0.707117), (33555,-0.335465), (33556,-0.520277), (33557,-0.392948), (33558,-0.531776), (33559,-0.511281), (33560,-0.440156), (33561,-0.618465), (33562,-0.664858), (33563,-0.416761), (33564,-0.417169), (33565,-0.602446), (33566,-0.590312), (33567,-0.786737), (33568,-0.519130), (33569,-0.636591), (33570,-0.714105), (33571,-0.477156), (33572,-0.315919), (33573,-0.496551), (33574,-0.555949), (33575,-0.631605), (33576,-0.629690), (33577,-0.789420), (33578,-0.457249), (33579,-0.577032), (33580,-0.582549), (33581,-0.751104), (33582,-0.814219), (33583,-0.998102), (33584,-0.706342), (33585,-0.828912), (33586,-0.487916), (33587,-0.645787), (33588,-0.495235), (33589,-0.636384), (33590,-0.615425), (33591,-0.771903), (33592,-0.467137), (33593,-0.612467), (33594,-0.671866), (33595,-0.436775), (33596,-0.420461), (33597,-0.594590), (33598,-0.622403), (33599,-0.813718), (33600,-0.567479), (33601,-0.724421), (33602,-0.756878), (33603,-0.499027), (33604,-0.345687), (33605,-0.508204), (33606,-0.551345), (33607,-0.620962), (33608,-0.467622), (33609,-0.606450), (33610,-0.688608), (33611,-0.456768), (33612,-0.439525), (33613,-0.591823), (33614,-0.641003), (33615,-0.811415), (33616,-0.539629), (33617,-0.680779), (33618,-0.741571), (33619,-0.545961), (33620,-0.400518), (33621,-0.522159), (33622,-0.577842), (33623,-0.659536), (33624,-0.469501), (33625,-0.609721), (33626,-0.632889), (33627,-0.421023), (33628,-0.415857), (33629,-0.565367), (33630,-0.607579), (33631,-0.787746), (33632,-0.508993), (33633,-0.684515), (33634,-0.740662), (33635,-0.492565), (33636,-0.342476), (33637,-0.513819), (33638,-0.530484), (33639,-0.608926), (33640,-0.553595), (33641,-0.702640), (33642,-0.372328), (33643,-0.502794), (33644,-0.482764), (33645,-0.657357), (33646,-0.722330), (33647,-0.877414), (33648,-0.605164), (33649,-0.755603), (33650,-0.419252), (33651,-0.568763), (33652,-0.435860), (33653,-0.583513), (33654,-0.540258), (33655,-0.695807), (33656,-0.587523), (33657,-0.726814), (33658,-0.409508), (33659,-0.521859), (33660,-0.520408), (33661,-0.649016), (33662,-0.726995), (33663,-0.901588), (33664,-0.694367), (33665,-0.879179), (33666,-0.912566), (33667,-0.676545), (33668,-0.509271), (33669,-0.677361), (33670,-0.721431), (33671,-0.777114), (33672,-0.745936), (33673,-0.894982), (33674,-0.576746), (33675,-0.720218), (33676,-0.705762), (33677,-0.874317), (33678,-0.953689), (33679,-1.100412), (33680,-0.790073), (33681,-0.969776), (33682,-0.631567), (33683,-0.801050), (33684,-0.649568), (33685,-0.813014), (33686,-0.797164), (33687,-0.940172), (33688,-0.929431), (33689,-0.666471), (33690,-0.811801), (33691,-0.482417), (33692,-0.640289), (33693,-0.610039), (33694,-0.769305), (33695,-0.844960), (33696,-1.001439), (33697,-0.742658), (33698,-0.889846), (33699,-0.566965), (33700,-0.709508), (33701,-0.581716), (33702,-0.701498), (33703,-0.676359), (33704,-1.085522), (33705,-0.825812), (33706,-0.562852), (33707,-0.602741), (33708,-0.747143), (33709,-0.722003), (33710,-0.937007), (33711,-1.000586), (33712,-1.169141), (33713,-0.879704), (33714,-0.641826), (33715,-0.712373), (33716,-0.862812), (33717,-0.681602), (33718,-0.772587), (33719,-0.857067), (33720,-1.016333), (33721,-0.733863), (33722,-0.887089), (33723,-0.505683), (33724,-0.683992), (33725,-0.664891), (33726,-0.800466), (33727,-0.887735), (33728,-1.039103), (33729,-0.775677), (33730,-0.913576), (33731,-0.584192), (33732,-0.725806), (33733,-0.589188), (33734,-0.761923), (33735,-0.727494), (33736,-1.013566), (33737,-0.733883), (33738,-0.507153), (33739,-0.527998), (33740,-0.697947), (33741,-0.694639), (33742,-0.890134), (33743,-0.929559), (33744,-1.114371), (33745,-0.843049), (33746,-0.562902), (33747,-0.603721), (33748,-0.813151), (33749,-0.660741), (33750,-0.743828), (33751,-0.822271), (33752,-0.991290), (33753,-0.690241), (33754,-0.831855), (33755,-0.507581), (33756,-0.643157), (33757,-0.608263), (33758,-0.762418), (33759,-0.849222), (33760,-0.983404), (33761,-0.676781), (33762,-0.842084), (33763,-0.514094), (33764,-0.653850), (33765,-0.533025), (33766,-0.681606), (33767,-0.675511), (33768,-0.879367), (33769,-0.608975), (33770,-0.734796), (33771,-0.407735), (33772,-0.554459), (33773,-0.543718), (33774,-0.695551), (33775,-0.762846), (33776,-0.900280), (33777,-0.653112), (33778,-0.781256), (33779,-0.448621), (33780,-0.626001), (33781,-0.445720), (33782,-0.591515), (33783,-0.553370), (33784,-0.776270), (33785,-0.521206), (33786,-0.650278), (33787,-0.330649), (33788,-0.479695), (33789,-0.450375), (33790,-0.586415), (33791,-0.659284), (33792,-0.819942), (33793,-0.547227), (33794,-0.683732), (33795,-0.356207), (33796,-0.517794), (33797,-0.355628), (33798,-0.487953), (33799,-0.467923), (33800,-0.800444), (33801,-0.540735), (33802,-0.711612), (33803,-0.365507), (33804,-0.515946), (33805,-0.502883), (33806,-0.675154), (33807,-0.762887), (33808,-0.890566), (33809,-0.606239), (33810,-0.737169), (33811,-0.393386), (33812,-0.568444), (33813,-0.439722), (33814,-0.583659), (33815,-0.545514), (33816,-0.591906), (33817,-0.753493), (33818,-0.794312), (33819,-0.563402), (33820,-0.548946), (33821,-0.718429), (33822,-0.796872), (33823,-0.947311), (33824,-0.690854), (33825,-0.813888), (33826,-0.857493), (33827,-0.653524), (33828,-0.479746), (33829,-0.655268), (33830,-0.733711), (33831,-0.801470), (33832,-0.532007), (33833,-0.685698), (33834,-0.730232), (33835,-0.481206), (33836,-0.488582), (33837,-0.635305), (33838,-0.664511), (33839,-0.863723), (33840,-0.613768), (33841,-0.770246), (33842,-0.801310), (33843,-0.575044), (33844,-0.410557), (33845,-0.575395), (33846,-0.652909), (33847,-0.716488), (33848,-0.530169), (33849,-0.648094), (33850,-0.696809), (33851,-0.441744), (33852,-0.444010), (33853,-0.593521), (33854,-0.647345), (33855,-0.864207), (33856,-0.551081), (33857,-0.726139), (33858,-0.754416), (33859,-0.514680), (33860,-0.387352), (33861,-0.572629), (33862,-0.623666), (33863,-0.712328), (33864,-0.525080), (33865,-0.685738), (33866,-0.732131), (33867,-0.447804), (33868,-0.426844), (33869,-0.596328), (33870,-0.628321), (33871,-0.813134), (33872,-0.563643), (33873,-0.749384), (33874,-0.782306), (33875,-0.552324), (33876,-0.396662), (33877,-0.514587), (33878,-0.547974), (33879,-0.659396), (33880,-0.552041), (33881,-0.745213), (33882,-0.789749), (33883,-0.546296), (33884,-0.510938), (33885,-0.719904), (33886,-0.785805), (33887,-0.919523), (33888,-0.629621), (33889,-0.805608), (33890,-0.858503), (33891,-0.607620), (33892,-0.459854), (33893,-0.614009), (33894,-0.657615), (33895,-0.722587), (33896,-0.680261), (33897,-0.817695), (33898,-0.452545), (33899,-0.602056), (33900,-0.608967), (33901,-0.756619), (33902,-0.842494), (33903,-0.995720), (33904,-0.696064), (33905,-0.856723), (33906,-0.481819), (33907,-0.649909), (33908,-0.487744), (33909,-0.622391), (33910,-0.593999), (33911,-0.770451), (33912,-0.519102), (33913,-0.686264), (33914,-0.706644), (33915,-0.474340), (33916,-0.459884), (33917,-0.634477), (33918,-0.691089), (33919,-0.893552), (33920,-0.725813), (33921,-0.870678), (33922,-0.967236), (33923,-0.720068), (33924,-0.550471), (33925,-0.727387), (33926,-0.774244), (33927,-0.822959), (33928,-0.656148), (33929,-0.833529), (33930,-0.900359), (33931,-0.635076), (33932,-0.603433), (33933,-0.747834), (33934,-0.789582), (33935,-0.986935), (33936,-0.679383), (33937,-0.846080), (33938,-0.899440), (33939,-0.642053), (33940,-0.496145), (33941,-0.630792), (33942,-0.727814), (33943,-0.796967), (33944,-0.961806), (33945,-0.670047), (33946,-0.839066), (33947,-0.471129), (33948,-0.633181), (33949,-0.639163), (33950,-0.740830), (33951,-0.837853), (33952,-0.991544), (33953,-0.714184), (33954,-0.872520), (33955,-0.528737), (33956,-0.647591), (33957,-0.521191), (33958,-0.676276), (33959,-0.633021), (33960,-1.058441), (33961,-0.808486), (33962,-0.545990), (33963,-0.581235), (33964,-0.755364), (33965,-0.737656), (33966,-0.909462), (33967,-0.977222), (33968,-1.126732), (33969,-0.852623), (33970,-0.608707), (33971,-0.677860), (33972,-0.837125), (33973,-0.655450), (33974,-0.765014), (33975,-0.818375), (33976,-0.978568), (33977,-0.700279), (33978,-0.852113), (33979,-0.506007), (33980,-0.679672), (33981,-0.673576), (33982,-0.811010), (33983,-0.877840), (33984,-1.016667), (33985,-0.746739), (33986,-0.899501), (33987,-0.550144), (33988,-0.694545), (33989,-0.578365), (33990,-0.744597), (33991,-0.714348), (33992,-0.909379), (33993,-0.629697), (33994,-0.797322), (33995,-0.458184), (33996,-0.649964), (33997,-0.628541), (33998,-0.759471), (33999,-0.839772), (34000,-0.998108), (34001,-0.703097), (34002,-0.832169), (34003,-0.490709), (34004,-0.673663), (34005,-0.535187), (34006,-0.654970), (34007,-0.624257), (34008,-0.908935), (34009,-0.673379), (34010,-0.801523), (34011,-0.470746), (34012,-0.614682), (34013,-0.578859), (34014,-0.757169), (34015,-0.823535), (34016,-0.985122), (34017,-0.724484), (34018,-0.889322), (34019,-0.528818), (34020,-0.690405), (34021,-0.553787), (34022,-0.698653), (34023,-0.700454), (34024,-0.845784), (34025,-0.572140), (34026,-0.706786), (34027,-0.374616), (34028,-0.540384), (34029,-0.549617), (34030,-0.703772), (34031,-0.750629), (34032,-0.909430), (34033,-0.663191), (34034,-0.811773), (34035,-0.466596), (34036,-0.633757), (34037,-0.468341), (34038,-0.615064), (34039,-0.576454), (34040,-0.835585), (34041,-0.591204), (34042,-0.730961), (34043,-0.393216), (34044,-0.539475), (34045,-0.493898), (34046,-0.682891), (34047,-0.804067), (34048,-0.943358), (34049,-0.646954), (34050,-0.840127), (34051,-0.478229), (34052,-0.604050), (34053,-0.463716), (34054,-0.606259), (34055,-0.576474), (34056,-0.897848), (34057,-0.628384), (34058,-0.755134), (34059,-0.408565), (34060,-0.562256), (34061,-0.550587), (34062,-0.701026), (34063,-0.777146), (34064,-0.941985), (34065,-0.666947), (34066,-0.838754), (34067,-0.496829), (34068,-0.670493), (34069,-0.513901), (34070,-0.696856), (34071,-0.675897), (34072,-0.588515), (34073,-0.745457), (34074,-0.801604), (34075,-0.566513), (34076,-0.566456), (34077,-0.720147), (34078,-0.768862), (34079,-0.925340), (34080,-0.623827), (34081,-0.787272), (34082,-0.898229), (34083,-0.658958), (34084,-0.470316), (34085,-0.634226), (34086,-0.665755), (34087,-0.755345), (34088,-0.516538), (34089,-0.675803), (34090,-0.730556), (34091,-0.499646), (34092,-0.479616), (34093,-0.646777), (34094,-0.673661), (34095,-0.860796), (34096,-0.593190), (34097,-0.731553), (34098,-0.780268), (34099,-0.527062), (34100,-0.368612), (34101,-0.526483), (34102,-0.591456), (34103,-0.682440), (34104,-0.573691), (34105,-0.716699), (34106,-0.787710), (34107,-0.559122), (34108,-0.492178), (34109,-0.657017), (34110,-0.693655), (34111,-0.904014), (34112,-0.638266), (34113,-0.779416), (34114,-0.842066), (34115,-0.632058), (34116,-0.500549), (34117,-0.652382), (34118,-0.717354), (34119,-0.758173), (34120,-0.609478), (34121,-0.749234), (34122,-0.791910), (34123,-0.551710), (34124,-0.523783), (34125,-0.680726), (34126,-0.763349), (34127,-0.929117), (34128,-0.651293), (34129,-0.790584), (34130,-0.849054), (34131,-0.622788), (34132,-0.483383), (34133,-0.665408), (34134,-0.662100), (34135,-0.762838), (34136,-0.592312), (34137,-0.716275), (34138,-0.758952), (34139,-0.520610), (34140,-0.551674), (34141,-0.692823), (34142,-0.735500), (34143,-0.925886), (34144,-0.636914), (34145,-0.776669), (34146,-0.853254), (34147,-0.632098), (34148,-0.461107), (34149,-0.598077), (34150,-0.646327), (34151,-0.701080), (34152,-0.676870), (34153,-0.809659), (34154,-0.457980), (34155,-0.608884), (34156,-0.605111), (34157,-0.750905), (34158,-0.844212), (34159,-0.998368), (34160,-0.730297), (34161,-0.884917), (34162,-0.560178), (34163,-0.714799), (34164,-0.569819), (34165,-0.757883), (34166,-0.696977), (34167,-0.852991), (34168,-0.589566), (34169,-0.726534), (34170,-0.762244), (34171,-0.488600), (34172,-0.463460), (34173,-0.621332), (34174,-0.670976), (34175,-0.852072), (34176,-0.975106), (34177,-0.671270), (34178,-0.824496), (34179,-0.526234), (34180,-0.685499), (34181,-0.547023), (34182,-0.710468), (34183,-0.667678), (34184,-1.029462), (34185,-0.728877), (34186,-0.497038), (34187,-0.542501), (34188,-0.717095), (34189,-0.702174), (34190,-0.918572), (34191,-0.969609), (34192,-1.142809), (34193,-0.838973), (34194,-0.623391), (34195,-0.666996), (34196,-0.788637), (34197,-0.637620), (34198,-0.712811), (34199,-0.791718), (34200,-0.898495), (34201,-0.628567), (34202,-0.774826), (34203,-0.404102), (34204,-0.527136), (34205,-0.554950), (34206,-0.685880), (34207,-0.779187), (34208,-0.910582), (34209,-0.623932), (34210,-0.780874), (34211,-0.477502), (34212,-0.594034), (34213,-0.434191), (34214,-0.584166), (34215,-0.615231), (34216,-1.033219), (34217,-0.778619), (34218,-0.530987), (34219,-0.582488), (34220,-0.739895), (34221,-0.756096), (34222,-0.911645), (34223,-0.951999), (34224,-1.134024), (34225,-0.846910), (34226,-0.611354), (34227,-0.681436), (34228,-0.799826), (34229,-0.645092), (34230,-0.748153), (34231,-0.773643), (34232,-0.966352), (34233,-0.700140), (34234,-0.872410), (34235,-0.553246), (34236,-0.674422), (34237,-0.703628), (34238,-0.829449), (34239,-0.915324), (34240,-1.052293), (34241,-0.772146), (34242,-0.923050), (34243,-0.583913), (34244,-0.689760), (34245,-0.528989), (34246,-0.673854), (34247,-0.685410), (34248,-1.012357), (34249,-0.708521), (34250,-0.469714), (34251,-0.524932), (34252,-0.667939), (34253,-0.619110), (34254,-0.820644), (34255,-0.911629), (34256,-1.056029), (34257,-0.754980), (34258,-0.485981), (34259,-0.576501), (34260,-0.722759), (34261,-0.601005), (34262,-0.654366), (34263,-0.696578), (34264,-0.892537), (34265,-0.622609), (34266,-0.783268), (34267,-0.444130), (34268,-0.588531), (34269,-0.584758), (34270,-0.755635), (34271,-0.834543), (34272,-0.966403), (34273,-0.726666), (34274,-0.862242), (34275,-0.487803), (34276,-0.662860), (34277,-0.488618), (34278,-0.659495), (34279,-0.622743), (34280,-0.675174), (34281,-0.831652), (34282,-0.545931), (34283,-0.321988), (34284,-0.373955), (34285,-0.542045), (34286,-0.540595), (34287,-0.699395), (34288,-0.767619), (34289,-0.935709), (34290,-0.646737), (34291,-0.410717), (34292,-0.467793), (34293,-0.618697), (34294,-0.478827), (34295,-0.541477), (34296,-0.745798), (34297,-0.477263), (34298,-0.623987), (34299,-0.260695), (34300,-0.438540), (34301,-0.422226), (34302,-0.545260), (34303,-0.663649), (34304,-0.773678), (34305,-0.519078), (34306,-0.643041), (34307,-0.321090), (34308,-0.453414), (34309,-0.327479), (34310,-0.460732), (34311,-0.416084), (34312,-0.631553), (34313,-0.797321), (34314,-0.523212), (34315,-0.294159), (34316,-0.348913), (34317,-0.527222), (34318,-0.515088), (34319,-0.671566), (34320,-0.720746), (34321,-0.881404), (34322,-0.611476), (34323,-0.381958), (34324,-0.430209), (34325,-0.590403), (34326,-0.438921), (34327,-0.499713), (34328,-0.539603), (34329,-0.685862), (34330,-0.716462), (34331,-0.476261), (34332,-0.475276), (34333,-0.628502), (34334,-0.695333), (34335,-0.860171), (34336,-0.558658), (34337,-0.729999), (34338,-0.790791), (34339,-0.556629), (34340,-0.386102), (34341,-0.534684), (34342,-0.599192), (34343,-0.675312), (34344,-0.792773), (34345,-0.500549), (34346,-0.655169), (34347,-0.314173), (34348,-0.472974), (34349,-0.450156), (34350,-0.546715), (34351,-0.665104), (34352,-0.816937), (34353,-0.556763), (34354,-0.693732), (34355,-0.323937), (34356,-0.471590), (34357,-0.346120), (34358,-0.486805), (34359,-0.463059), (34360,-0.379393), (34361,-0.551664), (34362,-0.613385), (34363,-0.364823), (34364,-0.352225), (34365,-0.528211), (34366,-0.578785), (34367,-0.738049), (34368,-0.478340), (34369,-0.628315), (34370,-0.692359), (34371,-0.448442), (34372,-0.303927), (34373,-0.443684), (34374,-0.505869), (34375,-0.585241), (34376,-0.743113), (34377,-0.460643), (34378,-0.589251), (34379,-0.252900), (34380,-0.413558), (34381,-0.429759), (34382,-0.573231), (34383,-0.590361), (34384,-0.759380), (34385,-0.506638), (34386,-0.663580), (34387,-0.328158), (34388,-0.513900), (34389,-0.317362), (34390,-0.491490), (34391,-0.443126), (34392,-0.459791), (34393,-0.587006), (34394,-0.661732), (34395,-0.431751), (34396,-0.411256), (34397,-0.570986), (34398,-0.635958), (34399,-0.796617), (34400,-0.511360), (34401,-0.685489), (34402,-0.723520), (34403,-0.503293), (34404,-0.343450), (34405,-0.505967), (34406,-0.530992), (34407,-0.604326), (34408,-0.885288), (34409,-0.571233), (34410,-0.367263), (34411,-0.409011), (34412,-0.574314), (34413,-0.583548), (34414,-0.753960), (34415,-0.790134), (34416,-0.955437), (34417,-0.684115), (34418,-0.451811), (34419,-0.510746), (34420,-0.673726), (34421,-0.479975), (34422,-0.566314), (34423,-0.609920), (34424,-0.785442), (34425,-0.520159), (34426,-0.645516), (34427,-0.317526), (34428,-0.464714), (34429,-0.493456), (34430,-0.656436), (34431,-0.728376), (34432,-1.007016), (34433,-0.733372), (34434,-0.852691), (34435,-0.527952), (34436,-0.687681), (34437,-0.518548), (34438,-0.691748), (34439,-0.690298), (34440,-0.921559), (34441,-0.656741), (34442,-0.816934), (34443,-0.455501), (34444,-0.626842), (34445,-0.594736), (34446,-0.768400), (34447,-0.813864), (34448,-0.990779), (34449,-0.702271), (34450,-0.890335), (34451,-0.549803), (34452,-0.697456), (34453,-0.523214), (34454,-0.692233), (34455,-0.641082), (34456,-0.896032), (34457,-0.631678), (34458,-0.753319), (34459,-0.444838), (34460,-0.584594), (34461,-0.560383), (34462,-0.724293), (34463,-0.794375), (34464,-0.962001), (34465,-0.659558), (34466,-0.795598), (34467,-0.460641), (34468,-0.589713), (34469,-0.466566), (34470,-0.614218), (34471,-0.572821), (34472,-0.930890), (34473,-1.071575), (34474,-0.392427), (34475,-0.554943), (34476,-0.584614), (34477,-0.769891), (34478,-0.775408), (34479,-0.931422), (34480,-0.978743), (34481,-1.123144), (34482,-0.475582), (34483,-0.638563), (34484,-0.715148), (34485,-0.860942), (34486,-0.628638), (34487,-0.767929), (34488,-0.936484), (34489,-0.634041), (34490,-0.814673), (34491,-0.471355), (34492,-0.619472), (34493,-0.609660), (34494,-0.790756), (34495,-0.868270), (34496,-1.039612), (34497,-0.703725), (34498,-0.855559), (34499,-0.550793), (34500,-0.750005), (34501,-0.586446), (34502,-0.733169), (34503,-0.692237), (34504,-0.792511), (34505,-0.978717), (34506,-0.682312), (34507,-0.436538), (34508,-0.479679), (34509,-0.631512), (34510,-0.585935), (34511,-0.786075), (34512,-0.836648), (34513,-0.967579), (34514,-0.726450), (34515,-0.475101), (34516,-0.533106), (34517,-0.711415), (34518,-0.579907), (34519,-0.649523), (34520,-0.920267), (34521,-0.636869), (34522,-0.778947), (34523,-0.425410), (34524,-0.586533), (34525,-0.609237), (34526,-0.784294), (34527,-0.852518), (34528,-0.993668), (34529,-0.708411), (34530,-0.883469), (34531,-0.542009), (34532,-0.710563), (34533,-0.531676), (34534,-0.664000), (34535,-0.621674), (34536,-0.721948), (34537,-0.894684), (34538,-0.600137), (34539,-0.321384), (34540,-0.351055), (34541,-0.501494), (34542,-0.498650), (34543,-0.699720), (34544,-0.730784), (34545,-0.851496), (34546,-0.580638), (34547,-0.378527), (34548,-0.426313), (34549,-0.598119), (34550,-0.411800), (34551,-0.495352), (34552,-0.790249), (34553,-0.524502), (34554,-0.649394), (34555,-0.285638), (34556,-0.456051), (34557,-0.478754), (34558,-0.599930), (34559,-0.713210), (34560,-0.865508), (34561,-0.577465), (34562,-0.722794), (34563,-0.393875), (34564,-0.582403), (34565,-0.428599), (34566,-0.579967), (34567,-0.532067), (34568,-0.753574), (34569,-0.905408), (34570,-0.635944), (34571,-0.382273), (34572,-0.419841), (34573,-0.557738), (34574,-0.543282), (34575,-0.744352), (34576,-0.812111), (34577,-0.977879), (34578,-0.706557), (34579,-0.466357), (34580,-0.504389), (34581,-0.640429), (34582,-0.483837), (34583,-0.552061), (34584,-0.834417), (34585,-0.581210), (34586,-0.759984), (34587,-0.407376), (34588,-0.576395), (34589,-0.553579), (34590,-0.710521), (34591,-0.778280), (34592,-0.931506), (34593,-0.669939), (34594,-0.812018), (34595,-0.449191), (34596,-0.626571), (34597,-0.517358), (34598,-0.652005), (34599,-0.596208), (34600,-0.765227), (34601,-0.479971), (34602,-0.642487), (34603,-0.268977), (34604,-0.387831), (34605,-0.396135), (34606,-0.543323), (34607,-0.676576), (34608,-0.812152), (34609,-0.547333), (34610,-0.690805), (34611,-0.335874), (34612,-0.499784), (34613,-0.360843), (34614,-0.506174), (34615,-0.468492), (34616,-0.806588), (34617,-0.514829), (34618,-0.701034), (34619,-0.367470), (34620,-0.509084), (34621,-0.531787), (34622,-0.682227), (34623,-0.755561), (34624,-0.924115), (34625,-0.645362), (34626,-0.791156), (34627,-0.478494), (34628,-0.629863), (34629,-0.459337), (34630,-0.593983), (34631,-0.557696), (34632,-0.799641), (34633,-0.549221), (34634,-0.690835), (34635,-0.335905), (34636,-0.503066), (34637,-0.469101), (34638,-0.612573), (34639,-0.737465), (34640,-0.874435), (34641,-0.600326), (34642,-0.749372), (34643,-0.435781), (34644,-0.573215), (34645,-0.431951), (34646,-0.588430), (34647,-0.577225), (34648,-0.798268), (34649,-0.517191), (34650,-0.670882), (34651,-0.308056), (34652,-0.454779), (34653,-0.445432), (34654,-0.577292), (34655,-0.684533), (34656,-0.829399), (34657,-0.575264), (34658,-0.720594), (34659,-0.370308), (34660,-0.500310), (34661,-0.341396), (34662,-0.493229), (34663,-0.479237), (34664,-0.811758), (34665,-0.509316), (34666,-0.315100), (34667,-0.367995), (34668,-0.519828), (34669,-0.514198), (34670,-0.717589), (34671,-0.786742), (34672,-0.913957), (34673,-0.628236), (34674,-0.398254), (34675,-0.432106), (34676,-0.611809), (34677,-0.438031), (34678,-0.534124), (34679,-0.602348), (34680,-0.781122), (34681,-0.483324), (34682,-0.631905), (34683,-0.267220), (34684,-0.442278), (34685,-0.417603), (34686,-0.595912), (34687,-0.681787), (34688,-0.952531), (34689,-0.631973), (34690,-0.786592), (34691,-0.470679), (34692,-0.638305), (34693,-0.463598), (34694,-0.614502), (34695,-0.551739), (34696,-0.822482), (34697,-0.593429), (34698,-0.727612), (34699,-0.394048), (34700,-0.542629), (34701,-0.533747), (34702,-0.715772), (34703,-0.774242), (34704,-0.946048), (34705,-0.676584), (34706,-0.825166), (34707,-0.473951), (34708,-0.625784), (34709,-0.469657), (34710,-0.624741), (34711,-0.575912), (34712,-0.916330), (34713,-0.666375), (34714,-0.826105), (34715,-0.470245), (34716,-0.615575), (34717,-0.637814), (34718,-0.799866), (34719,-0.893172), (34720,-1.026426), (34721,-0.736060), (34722,-0.876745), (34723,-0.546432), (34724,-0.706162), (34725,-0.583478), (34726,-0.766897), (34727,-0.693915), (34728,-0.778396), (34729,-0.948344), (34730,-0.714182), (34731,-0.469337), (34732,-0.508297), (34733,-0.637834), (34734,-0.627559), (34735,-0.844885), (34736,-0.890814), (34737,-1.031963), (34738,-0.767609), (34739,-0.530660), (34740,-0.597955), (34741,-0.762329), (34742,-0.592267), (34743,-0.645627), (34744,-0.939131), (34745,-0.648301), (34746,-0.805243), (34747,-0.465176), (34748,-0.596107), (34749,-0.571432), (34750,-0.707008), (34751,-0.774767), (34752,-0.955399), (34753,-0.684541), (34754,-0.814079), (34755,-0.477264), (34756,-0.666720), (34757,-0.496658), (34758,-0.682864), (34759,-0.670266), (34760,-0.767753), (34761,-0.926553), (34762,-0.663128), (34763,-0.421069), (34764,-0.490222), (34765,-0.646236), (34766,-0.628529), (34767,-0.756207), (34768,-0.816070), (34769,-0.971155), (34770,-0.689150), (34771,-0.470316), (34772,-0.497200), (34773,-0.666219), (34774,-0.540285), (34775,-0.601076), (34776,-0.980512), (34777,-0.698971), (34778,-0.842908), (34779,-0.523279), (34780,-0.688118), (34781,-0.683415), (34782,-0.810630), (34783,-0.887680), (34784,-1.033474), (34785,-0.781661), (34786,-0.949752), (34787,-0.590176), (34788,-0.771737), (34789,-0.630009), (34790,-0.734928), (34791,-0.701892), (34792,-0.789625), (34793,-0.931703), (34794,-0.647376), (34795,-0.441548), (34796,-0.480973), (34797,-0.662998), (34798,-0.631356), (34799,-0.806414), (34800,-0.858380), (34801,-0.967479), (34802,-0.713808), (34803,-0.469892), (34804,-0.539045), (34805,-0.703419), (34806,-0.542648), (34807,-0.615981), (34808,-0.792897), (34809,-0.513214), (34810,-0.659009), (34811,-0.290607), (34812,-0.453588), (34813,-0.461428), (34814,-0.641131), (34815,-0.685200), (34816,-1.089254), (34817,-0.806784), (34818,-0.961869), (34819,-0.633879), (34820,-0.792215), (34821,-0.652810), (34822,-0.806501), (34823,-0.775787), (34824,-0.957812), (34825,-1.119400), (34826,-0.842040), (34827,-0.604161), (34828,-0.619898), (34829,-0.803781), (34830,-0.792576), (34831,-0.955557), (34832,-1.033535), (34833,-1.193729), (34834,-0.888499), (34835,-0.665485), (34836,-0.745321), (34837,-0.881362), (34838,-0.726164), (34839,-0.771627), (34840,-0.595991), (34841,-0.726922), (34842,-0.803042), (34843,-0.959984), (34844,-0.573933), (34845,-0.700683), (34846,-0.753578), (34847,-0.906805), (34848,-0.651276), (34849,-0.793819), (34850,-0.882481), (34851,-1.038959), (34852,-0.485689), (34853,-0.644490), (34854,-0.699243), (34855,-0.823671), (34856,-1.022882), (34857,-0.768747), (34858,-0.918257), (34859,-0.540567), (34860,-0.738384), (34861,-0.726251), (34862,-0.885051), (34863,-0.941663), (34864,-1.106966), (34865,-0.855617), (34866,-1.002805), (34867,-0.626508), (34868,-0.795992), (34869,-0.656122), (34870,-0.796807), (34871,-0.791641), (34872,-0.721910), (34873,-0.883962), (34874,-0.952650), (34875,-0.720346), (34876,-0.724470), (34877,-0.873051), (34878,-0.918979), (34879,-1.067096), (34880,-0.778589), (34881,-0.934602), (34882,-0.971240), (34883,-0.763090), (34884,-0.646909), (34885,-0.786665), (34886,-0.843741), (34887,-0.926364), (34888,-1.061476), (34889,-0.766930), (34890,-0.903434), (34891,-0.561973), (34892,-0.696620), (34893,-0.689132), (34894,-0.870228), (34895,-0.935200), (34896,-1.089356), (34897,-0.820821), (34898,-0.972189), (34899,-0.659528), (34900,-0.821579), (34901,-0.681246), (34902,-0.828433), (34903,-0.808403), (34904,-0.622084), (34905,-0.740474), (34906,-0.780828), (34907,-0.949847), (34908,-0.552183), (34909,-0.694262), (34910,-0.761092), (34911,-0.914318), (34912,-0.662970), (34913,-0.796223), (34914,-0.848190), (34915,-1.002809), (34916,-0.462081), (34917,-0.609734), (34918,-0.696072), (34919,-0.863234), (34920,-1.023892), (34921,-0.752571), (34922,-0.890933), (34923,-0.527641), (34924,-0.697590), (34925,-0.695675), (34926,-0.844257), (34927,-0.915732), (34928,-1.097293), (34929,-0.783702), (34930,-0.923922), (34931,-0.588500), (34932,-0.747301), (34933,-0.596283), (34934,-0.715137), (34935,-0.663057), (34936,-0.983037), (34937,-0.748410), (34938,-0.896992), (34939,-0.533236), (34940,-0.680888), (34941,-0.691515), (34942,-0.839632), (34943,-0.914823), (34944,-1.358824), (34945,-1.068458), (34946,-0.862165), (34947,-0.918312), (34948,-1.060391), (34949,-0.911696), (34950,-0.965056), (34951,-1.007732), (34952,-1.192544), (34953,-0.920294), (34954,-0.697279), (34955,-0.719983), (34956,-0.869029), (34957,-0.862934), (34958,-1.026379), (34959,-1.086242), (34960,-1.256190), (34961,-0.983475), (34962,-0.737236), (34963,-0.783165), (34964,-0.947539), (34965,-0.773761), (34966,-0.869854), (34967,-0.916247), (34968,-1.254342), (34969,-0.978376), (34970,-0.744214), (34971,-0.811044), (34972,-0.949871), (34973,-0.934951), (34974,-1.147168), (34975,-1.200992), (34976,-1.343071), (34977,-1.049453), (34978,-0.792532), (34979,-0.860755), (34980,-0.988435), (34981,-0.864822), (34982,-0.915860), (34983,-0.952498), (34984,-1.058810), (34985,-1.197173), (34986,-0.557972), (34987,-0.736281), (34988,-0.779886), (34989,-0.949370), (34990,-0.953958), (34991,-1.066774), (34992,-1.136391), (34993,-1.291476), (34994,-0.621153), (34995,-0.788779), (34996,-0.886730), (34997,-1.004191), (34998,-0.766777), (34999,-0.931151), (35000,-1.328702), (35001,-1.045768), (35002,-0.780485), (35003,-0.841277), (35004,-0.983820), (35005,-0.981441), (35006,-1.179259), (35007,-1.240515), (35008,-1.377019), (35009,-1.120098), (35010,-0.874787), (35011,-0.909104), (35012,-1.072084), (35013,-0.928963), (35014,-1.008335), (35015,-1.065875), (35016,-1.056064), (35017,-1.190246), (35018,-0.499950), (35019,-0.689872), (35020,-0.758560), (35021,-0.863944), (35022,-0.888041), (35023,-1.092361), (35024,-1.132716), (35025,-1.299877), (35026,-0.604472), (35027,-0.767918), (35028,-0.798517), (35029,-0.940131), (35030,-0.739413), (35031,-0.896819), (35032,-1.305982), (35033,-1.023513), (35034,-0.771236), (35035,-0.787436), (35036,-0.975500), (35037,-0.955469), (35038,-1.142139), (35039,-1.193642), (35040,-1.340830), (35041,-1.044425), (35042,-0.812586), (35043,-0.884990), (35044,-1.030320), (35045,-0.882554), (35046,-0.953565), (35047,-1.022253), (35048,-1.063536), (35049,-1.237665), (35050,-0.531577), (35051,-0.673191), (35052,-0.737235), (35053,-0.889532), (35054,-0.916880), (35055,-1.084041), (35056,-1.147156), (35057,-1.354728), (35058,-0.622628), (35059,-0.772138), (35060,-0.841291), (35061,-0.981047), (35062,-0.751530), (35063,-0.894073), (35064,-0.944182), (35065,-0.664499), (35066,-0.841415), (35067,-0.478588), (35068,-0.637853), (35069,-0.658698), (35070,-0.797525), (35071,-0.835557), (35072,-0.959985), (35073,-0.701669), (35074,-0.855824), (35075,-0.506932), (35076,-0.655049), (35077,-0.486845), (35078,-0.676302), (35079,-0.662775), (35080,-0.900075), (35081,-1.100216), (35082,-0.797308), (35083,-0.558037), (35084,-0.595140), (35085,-0.752082), (35086,-0.735768), (35087,-0.905252), (35088,-0.930277), (35089,-1.092329), (35090,-0.849342), (35091,-0.567337), (35092,-0.666217), (35093,-0.783213), (35094,-0.643344), (35095,-0.700420), (35096,-0.975808), (35097,-0.731892), (35098,-0.853533), (35099,-0.491634), (35100,-0.677840), (35101,-0.665242), (35102,-0.828222), (35103,-0.866719), (35104,-1.022732), (35105,-0.756984), (35106,-0.883734), (35107,-0.543203), (35108,-0.697359), (35109,-0.569566), (35110,-0.702819), (35111,-0.692079), (35112,-1.129576), (35113,-0.822953), (35114,-0.598080), (35115,-0.664446), (35116,-0.842756), (35117,-0.823655), (35118,-0.986171), (35119,-0.990759), (35120,-1.148631), (35121,-0.898211), (35122,-0.693312), (35123,-0.736453), (35124,-0.886428), (35125,-0.698715), (35126,-0.780410), (35127,-0.863033), (35128,-0.991642), (35129,-0.698953), (35130,-0.813626), (35131,-0.469379), (35132,-0.645830), (35133,-0.623478), (35134,-0.746977), (35135,-0.845392), (35136,-1.001870), (35137,-0.714291), (35138,-0.895852), (35139,-0.553927), (35140,-0.689967), (35141,-0.565891), (35142,-0.687067), (35143,-0.659605), (35144,-0.909911), (35145,-0.641841), (35146,-0.787170), (35147,-0.461503), (35148,-0.624019), (35149,-0.588661), (35150,-0.761396), (35151,-0.840303), (35152,-0.981917), (35153,-0.696196), (35154,-0.838740), (35155,-0.538154), (35156,-0.659795), (35157,-0.525499), (35158,-0.673152), (35159,-0.642903), (35160,-0.884383), (35161,-0.595876), (35162,-0.724949), (35163,-0.417861), (35164,-0.607782), (35165,-0.576605), (35166,-0.715896), (35167,-0.780868), (35168,-0.954997), (35169,-0.698074), (35170,-0.863842), (35171,-0.524240), (35172,-0.638914), (35173,-0.538991), (35174,-0.654128), (35175,-0.650820), (35176,-1.017250), (35177,-0.763114), (35178,-0.483432), (35179,-0.524250), (35180,-0.709527), (35181,-0.684852), (35182,-0.858052), (35183,-0.897941), (35184,-1.062315), (35185,-0.777988), (35186,-0.553116), (35187,-0.627378), (35188,-0.761561), (35189,-0.615188), (35190,-0.701527), (35191,-0.741881), (35192,-1.127819), (35193,-0.844421), (35194,-0.594931), (35195,-0.644575), (35196,-0.790834), (35197,-0.770339), (35198,-0.988595), (35199,-1.053567), (35200,-0.996378), (35201,-1.149140), (35202,-0.845767), (35203,-0.990633), (35204,-0.829861), (35205,-0.971476), (35206,-0.952839), (35207,-1.096311), (35208,-1.247215), (35209,-0.981002), (35210,-0.772387), (35211,-0.816923), (35212,-0.939956), (35213,-0.955693), (35214,-1.115887), (35215,-1.162744), (35216,-1.324331), (35217,-1.068802), (35218,-0.843930), (35219,-0.848054), (35220,-1.004067), (35221,-0.847475), (35222,-0.920345), (35223,-1.000645), (35224,-1.287181), (35225,-0.982417), (35226,-0.726423), (35227,-0.781177), (35228,-0.936261), (35229,-0.908334), (35230,-1.121481), (35231,-1.170661), (35232,-1.305307), (35233,-1.032127), (35234,-0.807720), (35235,-0.863867), (35236,-1.003623), (35237,-0.840993), (35238,-0.908752), (35239,-0.959790), (35240,-1.169220), (35241,-0.876997), (35242,-0.648408), (35243,-0.695730), (35244,-0.848027), (35245,-0.819172), (35246,-0.976579), (35247,-1.018791), (35248,-1.236118), (35249,-0.964796), (35250,-0.735743), (35251,-0.751015), (35252,-0.919570), (35253,-0.738360), (35254,-0.867433), (35255,-0.896639), (35256,-1.308589), (35257,-1.031229), (35258,-0.775236), (35259,-0.832312), (35260,-0.983216), (35261,-0.945534), (35262,-1.099690), (35263,-1.222724), (35264,-1.376880), (35265,-1.073972), (35266,-0.822624), (35267,-0.890384), (35268,-1.054758), (35269,-0.899095), (35270,-0.951526), (35271,-1.024860), (35272,-1.209207), (35273,-0.946246), (35274,-0.692111), (35275,-0.720853), (35276,-0.881047), (35277,-0.892138), (35278,-1.087169), (35279,-1.148425), (35280,-1.272388), (35281,-1.001996), (35282,-0.784556), (35283,-0.846277), (35284,-0.996252), (35285,-0.868459), (35286,-0.906955), (35287,-0.979824), (35288,-1.277508), (35289,-0.994110), (35290,-0.764593), (35291,-0.804018), (35292,-0.944703), (35293,-0.941859), (35294,-1.128530), (35295,-1.173993), (35296,-1.346263), (35297,-1.046608), (35298,-0.809659), (35299,-0.870915), (35300,-1.011136), (35301,-0.845719), (35302,-0.918123), (35303,-0.995638), (35304,-1.109846), (35305,-0.833415), (35306,-0.602040), (35307,-0.647039), (35308,-0.824884), (35309,-0.799280), (35310,-0.992452), (35311,-1.049528), (35312,-1.223658), (35313,-0.980670), (35314,-0.705168), (35315,-0.755276), (35316,-0.893639), (35317,-0.763060), (35318,-0.839180), (35319,-0.908797), (35320,-0.970983), (35321,-0.691764), (35322,-0.835701), (35323,-0.497957), (35324,-0.632603), (35325,-0.646481), (35326,-0.780199), (35327,-0.831701), (35328,-0.947303), (35329,-0.704316), (35330,-0.873335), (35331,-0.526765), (35332,-0.682779), (35333,-0.549412), (35334,-0.717967), (35335,-0.725342), (35336,-0.988654), (35337,-0.708971), (35338,-0.856159), (35339,-0.512841), (35340,-0.710659), (35341,-0.684126), (35342,-0.824346), (35343,-0.903718), (35344,-1.077382), (35345,-0.774475), (35346,-0.920734), (35347,-0.603892), (35348,-0.775698), (35349,-0.606565), (35350,-0.768617), (35351,-0.711428), (35352,-0.667243), (35353,-0.814896), (35354,-0.869649), (35355,-0.621553), (35356,-0.631250), (35357,-0.815133), (35358,-0.881964), (35359,-1.038442), (35360,-0.753650), (35361,-0.905947), (35362,-0.954662), (35363,-0.719572), (35364,-0.557870), (35365,-0.736179), (35366,-0.757490), (35367,-0.787160), (35368,-0.758305), (35369,-0.912925), (35370,-0.566355), (35371,-0.705647), (35372,-0.718131), (35373,-0.872287), (35374,-0.933079), (35375,-1.078409), (35376,-0.812661), (35377,-0.978893), (35378,-0.618389), (35379,-0.769757), (35380,-0.628494), (35381,-0.766392), (35382,-0.714311), (35383,-0.882402), (35384,-0.603649), (35385,-0.782422), (35386,-0.800945), (35387,-0.578395), (35388,-0.577874), (35389,-0.720417), (35390,-0.771455), (35391,-0.941403), (35392,-0.669153), (35393,-0.842352), (35394,-0.881778), (35395,-0.676414), (35396,-0.511926), (35397,-0.692557), (35398,-0.737092), (35399,-0.788130), (35400,-0.604598), (35401,-0.763398), (35402,-0.813507), (35403,-0.579344), (35404,-0.567675), (35405,-0.751558), (35406,-0.800738), (35407,-0.958610), (35408,-0.671959), (35409,-0.824257), (35410,-0.877152), (35411,-0.621159), (35412,-0.479896), (35413,-0.646593), (35414,-0.702740), (35415,-0.772357), (35416,-0.603689), (35417,-0.770385), (35418,-0.799127), (35419,-0.567753), (35420,-0.548652), (35421,-0.710239), (35422,-0.771031), (35423,-0.950734), (35424,-0.655258), (35425,-0.804304), (35426,-0.841871), (35427,-0.622573), (35428,-0.491993), (35429,-0.644755), (35430,-0.717160), (35431,-0.768662), (35432,-1.034760), (35433,-0.724885), (35434,-0.509303), (35435,-0.558018), (35436,-0.682911), (35437,-0.676351), (35438,-0.870917), (35439,-0.948431), (35440,-1.101657), (35441,-0.821046), (35442,-0.601748), (35443,-0.639780), (35444,-0.760956), (35445,-0.612261), (35446,-0.687917), (35447,-0.756605), (35448,-0.857808), (35449,-0.996635), (35450,-0.670503), (35451,-0.821871), (35452,-0.795803), (35453,-0.954604), (35454,-1.043265), (35455,-1.190918), (35456,-1.287011), (35457,-1.006864), (35458,-0.775025), (35459,-0.849751), (35460,-0.970463), (35461,-0.850567), (35462,-0.925293), (35463,-0.960074), (35464,-1.225708), (35465,-0.896324), (35466,-0.662627), (35467,-0.706697), (35468,-0.872930), (35469,-0.877053), (35470,-1.030744), (35471,-1.118012), (35472,-1.281458), (35473,-0.988304), (35474,-0.720234), (35475,-0.770808), (35476,-0.963516), (35477,-0.815750), (35478,-0.900696), (35479,-0.944301), (35480,-1.057581), (35481,-1.216846), (35482,-0.511222), (35483,-0.666771), (35484,-0.750788), (35485,-0.909588), (35486,-0.949942), (35487,-1.097130), (35488,-1.172786), (35489,-1.304646), (35490,-0.641755), (35491,-0.784763), (35492,-0.837658), (35493,-0.982988), (35494,-0.775303), (35495,-0.910878), (35496,-1.232716), (35497,-0.983226), (35498,-0.722123), (35499,-0.832152), (35500,-0.910594), (35501,-1.084723), (35502,-1.057261), (35503,-1.230461), (35504,-1.279176), (35505,-1.019931), (35506,-0.728172), (35507,-0.930170), (35508,-0.975633), (35509,-1.053612), (35510,-0.875654), (35511,-1.029344), (35512,-1.107788), (35513,-1.248937), (35514,-0.573505), (35515,-0.720228), (35516,-0.774982), (35517,-0.946324), (35518,-0.938371), (35519,-1.106925), (35520,-1.158427), (35521,-1.327911), (35522,-0.651550), (35523,-0.772262), (35524,-0.841415), (35525,-0.994641), (35526,-0.781846), (35527,-0.907667), (35528,-0.989362), (35529,-1.149555), (35530,-0.473659), (35531,-0.618525), (35532,-0.714618), (35533,-0.855767), (35534,-0.884045), (35535,-1.038665), (35536,-1.097134), (35537,-1.267082), (35538,-0.557743), (35539,-0.702608), (35540,-0.762936), (35541,-0.915698), (35542,-0.701044), (35543,-0.832439), (35544,-1.045585), (35545,-1.205779), (35546,-0.560075), (35547,-0.701225), (35548,-0.774093), (35549,-0.887838), (35550,-0.897536), (35551,-1.111611), (35552,-1.147320), (35553,-1.320985), (35554,-0.628366), (35555,-0.807140), (35556,-0.846565), (35557,-1.016513), (35558,-0.786067), (35559,-0.944867), (35560,-0.997763), (35561,-1.163531), (35562,-0.482989), (35563,-0.619959), (35564,-0.673318), (35565,-0.814468), (35566,-0.852964), (35567,-0.980179), (35568,-1.030288), (35569,-1.202558), (35570,-0.524804), (35571,-0.680818), (35572,-0.741609), (35573,-0.895300), (35574,-0.662996), (35575,-0.818545), (35576,-0.992674), (35577,-1.133359), (35578,-0.502054), (35579,-0.652029), (35580,-0.708176), (35581,-0.846074), (35582,-0.846017), (35583,-0.995063), (35584,-1.083261), (35585,-1.212797), (35586,-0.507638), (35587,-0.677586), (35588,-0.708186), (35589,-0.874419), (35590,-0.649546), (35591,-0.828320), (35592,-1.055866), (35593,-1.203053), (35594,-0.533660), (35595,-0.669700), (35596,-0.756039), (35597,-0.861887), (35598,-0.873907), (35599,-1.057790), (35600,-1.094893), (35601,-1.257410), (35602,-0.579190), (35603,-0.719875), (35604,-0.806679), (35605,-0.956654), (35606,-0.710880), (35607,-0.853887), (35608,-1.002934), (35609,-0.726967), (35610,-0.878799), (35611,-0.530837), (35612,-0.658980), (35613,-0.647776), (35614,-0.814472), (35615,-0.884090), (35616,-1.035458), (35617,-0.797116), (35618,-0.904822), (35619,-0.569864), (35620,-0.736096), (35621,-0.589259), (35622,-0.749917), (35623,-0.697837), (35624,-1.028966), (35625,-0.779010), (35626,-0.533236), (35627,-0.564765), (35628,-0.728210), (35629,-0.732334), (35630,-0.871161), (35631,-0.937991), (35632,-1.119552), (35633,-0.822683), (35634,-0.571335), (35635,-0.623301), (35636,-0.794643), (35637,-0.642696), (35638,-0.740183), (35639,-0.805621), (35640,-1.124671), (35641,-0.835234), (35642,-0.589460), (35643,-0.634924), (35644,-0.822987), (35645,-0.836400), (35646,-1.003098), (35647,-1.027659), (35648,-1.199001), (35649,-0.920247), (35650,-0.693052), (35651,-0.714362), (35652,-0.856905), (35653,-0.735151), (35654,-0.820097), (35655,-0.872064), (35656,-1.122369), (35657,-0.855693), (35658,-0.607596), (35659,-0.627048), (35660,-0.790957), (35661,-0.757921), (35662,-0.927405), (35663,-0.965437), (35664,-1.136779), (35665,-0.881250), (35666,-0.658700), (35667,-0.688836), (35668,-0.856926), (35669,-0.720307), (35670,-0.801073), (35671,-0.838640), (35672,-0.902219), (35673,-0.626252), (35674,-0.778550), (35675,-0.430587), (35676,-0.578704), (35677,-0.570286), (35678,-0.757885), (35679,-0.828896), (35680,-0.977013), (35681,-0.712659), (35682,-0.881213), (35683,-0.538824), (35684,-0.679509), (35685,-0.527098), (35686,-0.688221), (35687,-0.644966), (35688,-1.172575), (35689,-0.448836), (35690,-0.585340), (35691,-0.641488), (35692,-0.791463), (35693,-0.825778), (35694,-1.020809), (35695,-1.096000), (35696,-1.239937), (35697,-0.556609), (35698,-0.719589), (35699,-0.760408), (35700,-0.920602), (35701,-0.705020), (35702,-0.860569), (35703,-0.907890), (35704,-1.115463), (35705,-0.812555), (35706,-0.557491), (35707,-0.593201), (35708,-0.765007), (35709,-0.745906), (35710,-0.923286), (35711,-0.987329), (35712,-1.294768), (35713,-1.431737), (35714,-0.751660), (35715,-0.896525), (35716,-0.954066), (35717,-1.114260), (35718,-0.909826), (35719,-1.042149), (35720,-1.196305), (35721,-1.359750), (35722,-0.669455), (35723,-0.819430), (35724,-0.848171), (35725,-1.008830), (35726,-1.016669), (35727,-1.163857), (35728,-1.231616), (35729,-1.385308), (35730,-0.714520), (35731,-0.862173), (35732,-0.926217), (35733,-1.079907), (35734,-0.857822), (35735,-1.050531), (35736,-1.053261), (35737,-1.212526), (35738,-0.943527), (35739,-0.687533), (35740,-0.730675), (35741,-0.902481), (35742,-0.907998), (35743,-1.085842), (35744,-1.131306), (35745,-1.275707), (35746,-0.996025), (35747,-0.766507), (35748,-0.831015), (35749,-0.965198), (35750,-0.796530), (35751,-0.860108), (35752,-1.182875), (35753,-1.218120), (35754,-0.974668), (35755,-0.654575), (35756,-0.819878), (35757,-0.908539), (35758,-1.065017), (35759,-1.061709), (35760,-1.253489), (35761,-1.333325), (35762,-1.096376), (35763,-0.800436), (35764,-0.939263), (35765,-0.986120), (35766,-1.094291), (35767,-0.908436), (35768,-1.246066), (35769,-1.299891), (35770,-1.062942), (35771,-0.759106), (35772,-0.952279), (35773,-0.972196), (35774,-1.146324), (35775,-1.124436), (35776,-1.310177), (35777,-1.367253), (35778,-1.121944), (35779,-0.854802), (35780,-0.968082), (35781,-1.015404), (35782,-1.085486), (35783,-0.934004), (35784,-1.117887), (35785,-1.171246), (35786,-0.960774), (35787,-0.656009), (35788,-0.841285), (35789,-0.890929), (35790,-1.085031), (35791,-1.061750), (35792,-1.223801), (35793,-1.261833), (35794,-1.013737), (35795,-0.701539), (35796,-0.871023), (35797,-0.945750), (35798,-1.029767), (35799,-0.853666), (35800,-1.034762), (35801,-1.126675), (35802,-1.247852), (35803,-0.581710), (35804,-0.717285), (35805,-0.762749), (35806,-0.921085), (35807,-0.953078), (35808,-1.096086), (35809,-1.161523), (35810,-1.291524), (35811,-0.608661), (35812,-0.791614), (35813,-0.851478), (35814,-0.976835), (35815,-0.777045), (35816,-0.910762), (35817,-0.953904), (35818,-1.112704), (35819,-0.457710), (35820,-0.616046), (35821,-0.642465), (35822,-0.821703), (35823,-0.803996), (35824,-0.978124), (35825,-1.051922), (35826,-1.201897), (35827,-0.535755), (35828,-0.713135), (35829,-0.745128), (35830,-0.889994), (35831,-0.621460), (35832,-0.815562), (35833,-0.884250), (35834,-1.034689), (35835,-0.369476), (35836,-0.551037), (35837,-0.593713), (35838,-0.758088), (35839,-0.815164), (35840,-0.934482), (35841,-0.976695), (35842,-1.145249), (35843,-0.466566), (35844,-0.610967), (35845,-0.669901), (35846,-0.810121), (35847,-0.594539), (35848,-0.884327), (35849,-0.925610), (35850,-1.124821), (35851,-0.437777), (35852,-0.576140), (35853,-0.629035), (35854,-0.797590), (35855,-0.776631), (35856,-0.921497), (35857,-0.982753), (35858,-1.134122), (35859,-0.482379), (35860,-0.630031), (35861,-0.715906), (35862,-0.846372), (35863,-0.612674), (35864,-0.951235), (35865,-1.139298), (35866,-0.834532), (35867,-0.583649), (35868,-0.639796), (35869,-0.822285), (35870,-0.814797), (35871,-1.007041), (35872,-1.047860), (35873,-1.197834), (35874,-0.933016), (35875,-0.695138), (35876,-0.756859), (35877,-0.905440), (35878,-0.755816), (35879,-0.796635), (35880,-0.881581), (35881,-1.033878), (35882,-0.742119), (35883,-0.508885), (35884,-0.581290), (35885,-0.727549), (35886,-0.710770), (35887,-0.901156), (35888,-0.932221), (35889,-1.096595), (35890,-0.832241), (35891,-0.571138), (35892,-0.610098), (35893,-0.785156), (35894,-0.651790), (35895,-0.713046), (35896,-0.878349), (35897,-1.047833), (35898,-0.769079), (35899,-0.489861), (35900,-0.549260), (35901,-0.706667), (35902,-0.694069), (35903,-0.853798), (35904,-0.911339), (35905,-1.051095), (35906,-0.762122), (35907,-0.547005), (35908,-0.620803), (35909,-0.761023), (35910,-0.622547), (35911,-0.686126), (35912,-0.807302), (35913,-0.971212), (35914,-0.705000), (35915,-0.468980), (35916,-0.532559), (35917,-0.709474), (35918,-0.688051), (35919,-0.856141), (35920,-0.916468), (35921,-1.065979), (35922,-0.804876), (35923,-0.582791), (35924,-0.640331), (35925,-0.787055), (35926,-0.639289), (35927,-0.688468), (35928,-0.942490), (35929,-1.078530), (35930,-0.797919), (35931,-0.568402), (35932,-0.616188), (35933,-0.770343), (35934,-0.752636), (35935,-0.915152), (35936,-0.963867), (35937,-1.130564), (35938,-0.850881), (35939,-0.624616), (35940,-0.676118), (35941,-0.846530), (35942,-0.695978), (35943,-0.750266), (35944,-1.000572), (35945,-1.119890), (35946,-0.497875), (35947,-0.637167), (35948,-0.689134), (35949,-0.865585), (35950,-0.876676), (35951,-1.039657), (35952,-1.092552), (35953,-1.247172), (35954,-0.566631), (35955,-0.724502), (35956,-0.790868), (35957,-0.915296), (35958,-0.710861), (35959,-0.860837), (35960,-1.066551), (35961,-1.255079), (35962,-0.591724), (35963,-0.736125), (35964,-0.775550), (35965,-0.931099), (35966,-0.938010), (35967,-1.092165), (35968,-1.213806), (35969,-1.372141), (35970,-1.082240), (35971,-0.869909), (35972,-0.899116), (35973,-1.068135), (35974,-0.883674), (35975,-0.985806), (35976,-1.263517), (35977,-1.411634), (35978,-0.739453), (35979,-0.912653), (35980,-0.926996), (35981,-1.094621), (35982,-1.105713), (35983,-1.274732), (35984,-1.328092), (35985,-1.490144), (35986,-0.818892), (35987,-0.994879), (35988,-1.023156), (35989,-1.178240), (35990,-0.969626), (35991,-1.096376), (35992,-1.126047), (35993,-1.258835), (35994,-0.988443), (35995,-0.735701), (35996,-0.815073), (35997,-0.979447), (35998,-1.002615), (35999,-1.188356), (36000,-1.211988), (36001,-1.375434), (36002,-1.071133), (36003,-0.843009), (36004,-0.870822), (36005,-1.045880), (36006,-0.890217), (36007,-0.981666), (36008,-1.277492), (36009,-1.324814), (36010,-1.066033), (36011,-0.781241), (36012,-0.924713), (36013,-1.008266), (36014,-1.174034), (36015,-1.179550), (36016,-1.346712), (36017,-1.360590), (36018,-1.138505), (36019,-0.869506), (36020,-1.000901), (36021,-1.039861), (36022,-1.128059), (36023,-0.995621), (36024,-1.186472), (36025,-1.237045), (36026,-1.411173), (36027,-0.698117), (36028,-0.842983), (36029,-0.913529), (36030,-1.067685), (36031,-1.078775), (36032,-1.212494), (36033,-1.259815), (36034,-1.374953), (36035,-0.710204), (36036,-0.881546), (36037,-0.924223), (36038,-1.062586), (36039,-0.814488), (36040,-1.167448), (36041,-1.258432), (36042,-0.995935), (36043,-0.719505), (36044,-0.871337), (36045,-0.918659), (36046,-1.119264), (36047,-1.116420), (36048,-1.268718), (36049,-1.312323), (36050,-1.081413), (36051,-0.787795), (36052,-0.962853), (36053,-0.983699), (36054,-1.053780), (36055,-0.893937), (36056,-1.085252), (36057,-1.134432), (36058,-1.297877), (36059,-0.623839), (36060,-0.819334), (36061,-0.879197), (36062,-1.044501), (36063,-1.032831), (36064,-1.199992), (36065,-1.251959), (36066,-1.398218), (36067,-0.710710), (36068,-0.829099), (36069,-0.917296), (36070,-1.064020), (36071,-0.863301), (36072,-1.012347), (36073,-1.076855), (36074,-1.254700), (36075,-0.579268), (36076,-0.697657), (36077,-0.786783), (36078,-0.907495), (36079,-0.897684), (36080,-1.054161), (36081,-1.108450), (36082,-1.265393), (36083,-0.606218), (36084,-0.746439), (36085,-0.812340), (36086,-0.981824), (36087,-0.706787), (36088,-0.903676), (36089,-0.977009), (36090,-1.099114), (36091,-0.446907), (36092,-0.654479), (36093,-0.705981), (36094,-0.832267), (36095,-0.858222), (36096,-1.016558), (36097,-1.023469), (36098,-1.189701), (36099,-0.520307), (36100,-0.696758), (36101,-0.716210), (36102,-0.854573), (36103,-0.639920), (36104,-0.961293), (36105,-1.005828), (36106,-1.129791), (36107,-0.487338), (36108,-0.635920), (36109,-0.682313), (36110,-0.845758), (36111,-0.844308), (36112,-0.959910), (36113,-1.041139), (36114,-1.219913), (36115,-0.525901), (36116,-0.656832), (36117,-0.729701), (36118,-0.887572), (36119,-0.673384), (36120,-1.049103), (36121,-1.251566), (36122,-0.937511), (36123,-0.678730), (36124,-0.736736), (36125,-0.882065), (36126,-0.878757), (36127,-1.059389), (36128,-1.084414), (36129,-1.239499), (36130,-0.969571), (36131,-0.731693), (36132,-0.805026), (36133,-0.960111), (36134,-0.807235), (36135,-0.921444), (36136,-0.963656), (36137,-1.104341), (36138,-0.855780), (36139,-0.620224), (36140,-0.691235), (36141,-0.813805), (36142,-0.779840), (36143,-0.958614), (36144,-1.006864), (36145,-1.174954), (36146,-0.895272), (36147,-0.665290), (36148,-0.713077), (36149,-0.815673), (36150,-0.691132), (36151,-0.765394), (36152,-0.937665), (36153,-1.095536), (36154,-0.855336), (36155,-0.618387), (36156,-0.664780), (36157,-0.820328), (36158,-0.838851), (36159,-0.993006), (36160,-1.031038), (36161,-1.174046), (36162,-0.885073), (36163,-0.666704), (36164,-0.746076), (36165,-0.904877), (36166,-0.738530), (36167,-0.802574), (36168,-0.964625), (36169,-1.124819), (36170,-0.853498), (36171,-0.638380), (36172,-0.666658), (36173,-0.851005), (36174,-0.830511), (36175,-1.012536), (36176,-1.044529), (36177,-1.212619), (36178,-0.919466), (36179,-0.683446), (36180,-0.715440), (36181,-0.884459), (36182,-0.743660), (36183,-0.776583), (36184,-1.042681), (36185,-1.194049), (36186,-0.902290), (36187,-0.656981), (36188,-0.731242), (36189,-0.873321), (36190,-0.850504), (36191,-1.011627), (36192,-1.071490), (36193,-1.260947), (36194,-1.016101), (36195,-0.755463), (36196,-0.759122), (36197,-0.943934), (36198,-0.826825), (36199,-0.906661), (36200,-1.136529), (36201,-1.273034), (36202,-0.601318), (36203,-0.735500), (36204,-0.781893), (36205,-0.929545), (36206,-0.940172), (36207,-1.117088), (36208,-1.175557), (36209,-1.308810), (36210,-0.658925), (36211,-0.787998), (36212,-0.873408), (36213,-0.989940), (36214,-0.745094), (36215,-0.932228), (36216,-1.018104), (36217,-1.175046), (36218,-0.890254), (36219,-0.638441), (36220,-0.702949), (36221,-0.843634), (36222,-0.838468), (36223,-1.001449), (36224,-1.176971), (36225,-1.351564), (36226,-1.058411), (36227,-0.865125), (36228,-0.885505), (36229,-1.026655), (36230,-0.880282), (36231,-0.945255), (36232,-1.102197), (36233,-1.284687), (36234,-0.970167), (36235,-0.745295), (36236,-0.810268), (36237,-0.990899), (36238,-0.971798), (36239,-1.139888), (36240,-1.181172), (36241,-1.354836), (36242,-1.053787), (36243,-0.804296), (36244,-0.881345), (36245,-1.045720), (36246,-0.870548), (36247,-0.913690), (36248,-1.144951), (36249,-1.328834), (36250,-1.075628), (36251,-0.806628), (36252,-0.858595), (36253,-1.022040), (36254,-1.058679), (36255,-1.242562), (36256,-1.256904), (36257,-1.409202), (36258,-1.122087), (36259,-0.853553), (36260,-0.942679), (36261,-1.095441), (36262,-0.961145), (36263,-1.030763), (36264,-1.115243), (36265,-1.167210), (36266,-1.319972), (36267,-0.643611), (36268,-0.777793), (36269,-0.840908), (36270,-0.967194), (36271,-0.992684), (36272,-1.130582), (36273,-1.192767), (36274,-1.345530), (36275,-0.685426), (36276,-0.855374), (36277,-0.899445), (36278,-0.984855), (36279,-0.780420), (36280,-1.138489), (36281,-1.187668), (36282,-1.333463), (36283,-0.684042), (36284,-0.860029), (36285,-0.907816), (36286,-1.059184), (36287,-1.081423), (36288,-1.223966), (36289,-1.292654), (36290,-1.434733), (36291,-0.791351), (36292,-0.912527), (36293,-0.972855), (36294,-1.164634), (36295,-0.943943), (36296,-1.129683), (36297,-1.178399), (36298,-1.325122), (36299,-0.654335), (36300,-0.787124), (36301,-0.850239), (36302,-1.011826), (36303,-1.012234), (36304,-1.157099), (36305,-1.221142), (36306,-1.376226), (36307,-0.698473), (36308,-0.867027), (36309,-0.913884), (36310,-1.032738), (36311,-0.829697), (36312,-1.286703), (36313,-1.315909), (36314,-1.456130), (36315,-0.793239), (36316,-0.980374), (36317,-1.028160), (36318,-1.199038), (36319,-1.192013), (36320,-1.328517), (36321,-1.404174), (36322,-1.547646), (36323,-0.890329), (36324,-1.048200), (36325,-1.064401), (36326,-1.191151), (36327,-0.976498), (36328,-1.129724), (36329,-1.157072), (36330,-1.349781), (36331,-0.689678), (36332,-0.828040), (36333,-0.871181), (36334,-0.962630), (36335,-1.042931), (36336,-1.181758), (36337,-1.233724), (36338,-1.381377), (36339,-0.699442), (36340,-0.836875), (36341,-0.886055), (36342,-1.019308), (36343,-0.800010), (36344,-0.912361), (36345,-0.950857), (36346,-1.097581), (36347,-0.807215), (36348,-0.560047), (36349,-0.609227), (36350,-0.767563), (36351,-0.746603), (36352,-0.952782), (36353,-1.008465), (36354,-1.138466), (36355,-0.882473), (36356,-0.618119), (36357,-0.661724), (36358,-0.807983), (36359,-0.644889), (36360,-0.882654), (36361,-0.940658), (36362,-1.105033), (36363,-0.843466), (36364,-0.577718), (36365,-0.632007), (36366,-0.780589), (36367,-0.815369), (36368,-0.982530), (36369,-1.021026), (36370,-1.183078), (36371,-0.934981), (36372,-0.688278), (36373,-0.733277), (36374,-0.893006), (36375,-0.721551), (36376,-0.911473), (36377,-1.062376), (36378,-0.820782), (36379,-0.954965), (36380,-0.597711), (36381,-0.739790), (36382,-0.742056), (36383,-0.911075), (36384,-0.983479), (36385,-1.138099), (36386,-0.830547), (36387,-0.991670), (36388,-0.650210), (36389,-0.788108), (36390,-0.651954), (36391,-0.811683), (36392,-1.061989), (36393,-1.206390), (36394,-0.947610), (36395,-0.672572), (36396,-0.736151), (36397,-0.907493), (36398,-0.889785), (36399,-1.017929), (36400,-1.077328), (36401,-1.245418), (36402,-0.949943), (36403,-0.706955), (36404,-0.744987), (36405,-0.904252), (36406,-0.761130), (36407,-0.890203), (36408,-0.916158), (36409,-1.028045), (36410,-0.768335), (36411,-0.923884), (36412,-0.574992), (36413,-0.725432), (36414,-0.694718), (36415,-0.833545), (36416,-0.932426), (36417,-1.094942), (36418,-0.840342), (36419,-0.989853), (36420,-0.668830), (36421,-0.828559), (36422,-0.665000), (36423,-0.845168), (36424,-0.916643), (36425,-1.045716), (36426,-0.756743), (36427,-0.902538), (36428,-0.550394), (36429,-0.699440), (36430,-0.691022), (36431,-0.848429), (36432,-0.931517), (36433,-1.072202), (36434,-0.791126), (36435,-0.981047), (36436,-0.641910), (36437,-0.780737), (36438,-0.624610), (36439,-0.796416), (36440,-0.847454), (36441,-1.015543), (36442,-0.735396), (36443,-0.862611), (36444,-0.525796), (36445,-0.687848), (36446,-0.708693), (36447,-0.870281), (36448,-0.926892), (36449,-1.096840), (36450,-0.789753), (36451,-0.929973), (36452,-0.589907), (36453,-0.779363), (36454,-0.659003), (36455,-0.800616), (36456,-0.980784), (36457,-1.131223), (36458,-0.852934), (36459,-0.587186), (36460,-0.626147), (36461,-0.801669), (36462,-0.789535), (36463,-0.992927), (36464,-1.042571), (36465,-1.212984), (36466,-0.957456), (36467,-0.674986), (36468,-0.750642), (36469,-0.913158), (36470,-0.758889), (36471,-0.818752), (36472,-1.058839), (36473,-1.218104), (36474,-0.917519), (36475,-0.698221), (36476,-0.741362), (36477,-0.882047), (36478,-0.818819), (36479,-0.993412), (36480,-1.156393), (36481,-1.216720), (36482,-1.418254), (36483,-0.720062), (36484,-0.882114), (36485,-0.916430), (36486,-1.051076), (36487,-0.820166), (36488,-1.210285), (36489,-1.309165), (36490,-1.025302), (36491,-0.783708), (36492,-0.939257), (36493,-0.939664), (36494,-1.125406), (36495,-1.097944), (36496,-1.279040), (36497,-1.350515), (36498,-1.104741), (36499,-0.819484), (36500,-0.949951), (36501,-1.025142), (36502,-1.106372), (36503,-0.953496), (36504,-1.101149), (36505,-1.151257), (36506,-1.323992), (36507,-0.640664), (36508,-0.830586), (36509,-0.891842), (36510,-1.019057), (36511,-1.017142), (36512,-1.143428), (36513,-1.207471), (36514,-1.405289), (36515,-0.716387), (36516,-0.834312), (36517,-0.893710), (36518,-1.012564), (36519,-0.770505), (36520,-1.162018), (36521,-1.228848), (36522,-0.995615), (36523,-0.725222), (36524,-0.871946), (36525,-0.896507), (36526,-1.128698), (36527,-1.093340), (36528,-1.259572), (36529,-1.336621), (36530,-1.025817), (36531,-0.793049), (36532,-0.930018), (36533,-0.956438), (36534,-1.013978), (36535,-0.865282), (36536,-1.064029), (36537,-1.128537), (36538,-1.304989), (36539,-0.635130), (36540,-0.800434), (36541,-0.843575), (36542,-1.015846), (36543,-1.018112), (36544,-1.195492), (36545,-1.254890), (36546,-1.377924), (36547,-0.722002), (36548,-0.897988), (36549,-0.938807), (36550,-1.095749), (36551,-0.834182), (36552,-1.154626), (36553,-1.223779), (36554,-0.964070), (36555,-0.678349), (36556,-0.862232), (36557,-0.919308), (36558,-1.094366), (36559,-1.096631), (36560,-1.253574), (36561,-1.309721), (36562,-1.066733), (36563,-0.777761), (36564,-0.941206), (36565,-1.009430), (36566,-1.038172), (36567,-0.886690), (36568,-1.062212), (36569,-1.096064), (36570,-1.279947), (36571,-0.602192), (36572,-0.770283), (36573,-0.847796), (36574,-0.973153), (36575,-1.021403), (36576,-1.173701), (36577,-1.223345), (36578,-1.349166), (36579,-0.684418), (36580,-0.860869), (36581,-0.927699), (36582,-1.096254), (36583,-0.851873), (36584,-0.880151), (36585,-1.041273), (36586,-1.083486), (36587,-0.841427), (36588,-0.567783), (36589,-0.688495), (36590,-0.759041), (36591,-0.933634), (36592,-0.926146), (36593,-1.098881), (36594,-1.184756), (36595,-0.870701), (36596,-0.593805), (36597,-0.800913), (36598,-0.832442), (36599,-0.897878), (36600,-0.899679), (36601,-0.976264), (36602,-1.084899), (36603,-0.448950), (36604,-0.614253), (36605,-0.637421), (36606,-0.783679), (36607,-0.820318), (36608,-0.944281), (36609,-0.996712), (36610,-1.124856), (36611,-0.455927), (36612,-0.643062), (36613,-0.677377), (36614,-0.825030), (36615,-0.587617), (36616,-0.803549), (36617,-0.931229), (36618,-0.994808), (36619,-0.757859), (36620,-0.480499), (36621,-0.631867), (36622,-0.718671), (36623,-0.887690), (36624,-0.874163), (36625,-1.011132), (36626,-1.078892), (36627,-0.827543), (36628,-0.516275), (36629,-0.671359), (36630,-0.729829), (36631,-0.829638), (36632,-0.961498), (36633,-1.131446), (36634,-0.839222), (36635,-0.582300), (36636,-0.660278), (36637,-0.795389), (36638,-0.776753), (36639,-0.991292), (36640,-1.051155), (36641,-1.217853), (36642,-0.901475), (36643,-0.638050), (36644,-0.699306), (36645,-0.864609), (36646,-0.713592), (36647,-0.780422), (36648,-0.894166), (36649,-0.937772), (36650,-1.132339), (36651,-0.434611), (36652,-0.599450), (36653,-0.666280), (36654,-0.792566), (36655,-0.804586), (36656,-0.972212), (36657,-1.011637), (36658,-1.158825), (36659,-0.503367), (36660,-0.646839), (36661,-0.744790), (36662,-0.868753), (36663,-0.660138), (36664,-0.930882), (36665,-1.080392), (36666,-0.779808), (36667,-0.537285), (36668,-0.569278), (36669,-0.722040), (36670,-0.691791), (36671,-0.867313), (36672,-0.971303), (36673,-1.112452), (36674,-0.845312), (36675,-0.539153), (36676,-0.604590), (36677,-0.745275), (36678,-0.579858), (36679,-0.648547), (36680,-0.832894), (36681,-0.873712), (36682,-1.017649), (36683,-0.371480), (36684,-0.537248), (36685,-0.603614), (36686,-0.745693), (36687,-0.725198), (36688,-0.859845), (36689,-0.930856), (36690,-1.092443), (36691,-0.440236), (36692,-0.613900), (36693,-0.671440), (36694,-0.829312), (36695,-0.620232), (36696,-0.957863), (36697,-1.115734), (36698,-0.801679), (36699,-0.568911), (36700,-0.625523), (36701,-0.738802), (36702,-0.750358), (36703,-0.933312), (36704,-0.967628), (36705,-1.137576), (36706,-0.850461), (36707,-0.610261), (36708,-0.675698), (36709,-0.800590), (36710,-0.669082), (36711,-0.751241), (36712,-0.992256), (36713,-1.042829), (36714,-0.817028), (36715,-0.561500), (36716,-0.717977), (36717,-0.771337), (36718,-0.942214), (36719,-0.927294), (36720,-1.066121), (36721,-1.143635), (36722,-0.896931), (36723,-0.591701), (36724,-0.754682), (36725,-0.795501), (36726,-0.867441), (36727,-0.712243), (36728,-0.946292), (36729,-0.986181), (36730,-1.178425), (36731,-0.476052), (36732,-0.631601), (36733,-0.678923), (36734,-0.836330), (36735,-0.855317), (36736,-0.826462), (36737,-0.883074), (36738,-0.640551), (36739,-0.363191), (36740,-0.505734), (36741,-0.555378), (36742,-0.644969), (36743,-0.451682), (36744,-0.750759), (36745,-0.808300), (36746,-0.588537), (36747,-0.260547), (36748,-0.424921), (36749,-0.466205), (36750,-0.688641), (36751,-0.650496), (36752,-0.816263), (36753,-0.871481), (36754,-0.581580), (36755,-0.303291), (36756,-0.468594), (36757,-0.551682), (36758,-0.581353), (36759,-0.452631), (36760,-0.719194), (36761,-0.787883), (36762,-0.576016), (36763,-0.290760), (36764,-0.419368), (36765,-0.486198), (36766,-0.650573), (36767,-0.622181), (36768,-0.771692), (36769,-0.830626), (36770,-0.584387), (36771,-0.326536), (36772,-0.455144), (36773,-0.499214), (36774,-0.588341), (36775,-0.423853), (36776,-0.702492), (36777,-0.491555), (36778,-0.521226), (36779,-0.675381), (36780,-0.428678), (36781,-0.617670), (36782,-0.659883), (36783,-0.847482), (36784,-0.859967), (36785,-0.618373), (36786,-0.653617), (36787,-0.813811), (36788,-0.527625), (36789,-0.604675), (36790,-0.645958), (36791,-0.803830), (36792,-0.727596), (36793,-0.852952), (36794,-0.504060), (36795,-0.644281), (36796,-0.328368), (36797,-0.515038), (36798,-0.614847), (36799,-0.751816), (36800,-0.743863), (36801,-0.903592), (36802,-0.569564), (36803,-0.717681), (36804,-0.438463), (36805,-0.601444), (36806,-0.551686), (36807,-0.732782), (36808,-0.628214), (36809,-0.763325), (36810,-0.423723), (36811,-0.584381), (36812,-0.293086), (36813,-0.454209), (36814,-0.546122), (36815,-0.685878), (36816,-0.692325), (36817,-0.845551), (36818,-0.513845), (36819,-0.627589), (36820,-0.360913), (36821,-0.549905), (36822,-0.514546), (36823,-0.664522), (36824,-0.683045), (36825,-0.812117), (36826,-0.453471), (36827,-0.599265), (36828,-0.322834), (36829,-0.485815), (36830,-0.568438), (36831,-0.732813), (36832,-0.713711), (36833,-0.846036), (36834,-0.539412), (36835,-0.668950), (36836,-0.377190), (36837,-0.541100), (36838,-0.513174), (36839,-0.662684), (36840,-0.529782), (36841,-0.663035), (36842,-0.330400), (36843,-0.525895), (36844,-0.251322), (36845,-0.428703), (36846,-0.495533), (36847,-0.609742), (36848,-0.642199), (36849,-0.741080), (36850,-0.426560), (36851,-0.565388), (36852,-0.288028), (36853,-0.422674), (36854,-0.453274), (36855,-0.600927), (36856,-0.580896), (36857,-0.698357), (36858,-0.364793), (36859,-0.514768), (36860,-0.239731), (36861,-0.413859), (36862,-0.479760), (36863,-0.641812), (36864,-0.616673), (36865,-0.783834), (36866,-0.444696), (36867,-0.580272), (36868,-0.308950), (36869,-0.440345), (36870,-0.379439), (36871,-0.539169), (36872,-0.554440), (36873,-0.710454), (36874,-0.385716), (36875,-0.538478), (36876,-0.284807), (36877,-0.398551), (36878,-0.511831), (36879,-0.647407), (36880,-0.653388), (36881,-0.795467), (36882,-0.470264), (36883,-0.587724), (36884,-0.393973), (36885,-0.505395), (36886,-0.465391), (36887,-0.646952), (36888,-0.671049), (36889,-0.725802), (36890,-0.487925), (36891,-0.228680), (36892,-0.390731), (36893,-0.403216), (36894,-0.615433), (36895,-0.620021), (36896,-0.769996), (36897,-0.801061), (36898,-0.592446), (36899,-0.335059), (36900,-0.496182), (36901,-0.566728), (36902,-0.615444), (36903,-0.460710), (36904,-0.650167), (36905,-0.681231), (36906,-0.487481), (36907,-0.191076), (36908,-0.362882), (36909,-0.421352), (36910,-0.599196), (36911,-0.536433), (36912,-0.660396), (36913,-0.731407), (36914,-0.525579), (36915,-0.245432), (36916,-0.388904), (36917,-0.446445), (36918,-0.504450), (36919,-0.327885), (36920,-0.718003), (36921,-0.776938), (36922,-0.550672), (36923,-0.252410), (36924,-0.401455), (36925,-0.409295), (36926,-0.641021), (36927,-0.632604), (36928,-0.809983), (36929,-0.819681), (36930,-0.578087), (36931,-0.320701), (36932,-0.437232), (36933,-0.476657), (36934,-0.556493), (36935,-0.413372), (36936,-0.654853), (36937,-0.714716), (36938,-0.481947), (36939,-0.189723), (36940,-0.356884), (36941,-0.407458), (36942,-0.581122), (36943,-0.565272), (36944,-0.728717), (36945,-0.789974), (36946,-0.569746), (36947,-0.290064), (36948,-0.420066), (36949,-0.465065), (36950,-0.553262), (36951,-0.389239), (36952,-0.659982), (36953,-0.704517), (36954,-0.482431), (36955,-0.204143), (36956,-0.352260), (36957,-0.419554), (36958,-0.560240), (36959,-0.564363), (36960,-0.714338), (36961,-0.741222), (36962,-0.547007), (36963,-0.291942), (36964,-0.421944), (36965,-0.446506), (36966,-0.512871), (36967,-0.300540), (36968,-0.681369), (36969,-0.318078), (36970,-0.455511), (36971,-0.206950), (36972,-0.368073), (36973,-0.455341), (36974,-0.585807), (36975,-0.640561), (36976,-0.778459), (36977,-0.421205), (36978,-0.597657), (36979,-0.328658), (36980,-0.438222), (36981,-0.431662), (36982,-0.563986), (36983,-0.428761), (36984,-0.597316), (36985,-0.638599), (36986,-0.429055), (36987,-0.171669), (36988,-0.330933), (36989,-0.382900), (36990,-0.555171), (36991,-0.524922), (36992,-0.715308), (36993,-0.904300), (36994,-0.333844), (36995,-0.510295), (36996,-0.568765), (36997,-0.701089), (36998,-0.336404), (36999,-0.484521), (37000,-0.627528), (37001,-0.705507), (37002,-0.457410), (37003,-0.401614), (37004,-0.551124), (37005,-0.621206), (37006,-0.794406), (37007,-0.504040), (37008,-0.649835), (37009,-0.696692), (37010,-0.476464), (37011,-0.350065), (37012,-0.523265), (37013,-0.589630), (37014,-0.658319), (37015,-0.364237), (37016,-0.687933), (37017,-0.732468), (37018,-0.495055), (37019,-0.455980), (37020,-0.638934), (37021,-0.700191), (37022,-0.888719), (37023,-0.614145), (37024,-0.804532), (37025,-0.854640), (37026,-0.600040), (37027,-0.456455), (37028,-0.640338), (37029,-0.641674), (37030,-0.674132), (37031,-0.447866), (37032,-0.638253), (37033,-0.700902), (37034,-0.412859), (37035,-0.382610), (37036,-0.562777), (37037,-0.646794), (37038,-0.822780), (37039,-0.607198), (37040,-0.729303), (37041,-0.768264), (37042,-0.541534), (37043,-0.368686), (37044,-0.544207), (37045,-0.593851), (37046,-0.678333), (37047,-0.389825), (37048,-0.673110), (37049,-0.710212), (37050,-0.465367), (37051,-0.483426), (37052,-0.623182), (37053,-0.704876), (37054,-0.875289), (37055,-0.590032), (37056,-0.733969), (37057,-0.791509), (37058,-0.554096), (37059,-0.380318), (37060,-0.575814), (37061,-0.617096), (37062,-0.695540), (37063,-0.387058), (37064,-0.563974), (37065,-0.634985), (37066,-0.385959), (37067,-0.418881), (37068,-0.569321), (37069,-0.598991), (37070,-0.766617), (37071,-0.496224), (37072,-0.646664), (37073,-0.683767), (37074,-0.430096), (37075,-0.294871), (37076,-0.437879), (37077,-0.469872), (37078,-0.564108), (37079,-0.277922), (37080,-0.682905), (37081,-0.763206), (37082,-0.515109), (37083,-0.514123), (37084,-0.678032), (37085,-0.731393), (37086,-0.890193), (37087,-0.608653), (37088,-0.769776), (37089,-0.836606), (37090,-0.601979), (37091,-0.440743), (37092,-0.609297), (37093,-0.671019), (37094,-0.738778), (37095,-0.455844), (37096,-0.649017), (37097,-0.638277), (37098,-0.391109), (37099,-0.389659), (37100,-0.584225), (37101,-0.635727), (37102,-0.806140), (37103,-0.514380), (37104,-0.655530), (37105,-0.722825), (37106,-0.488198), (37107,-0.344148), (37108,-0.504807), (37109,-0.559560), (37110,-0.614778), (37111,-0.298401), (37112,-0.521301), (37113,-0.582558), (37114,-0.347466), (37115,-0.344159), (37116,-0.518287), (37117,-0.544707), (37118,-0.742989), (37119,-0.445191), (37120,-0.662053), (37121,-0.681970), (37122,-0.473819), (37123,-0.296326), (37124,-0.465809), (37125,-0.522421), (37126,-0.616192), (37127,-0.299814), (37128,-0.592389), (37129,-0.652717), (37130,-0.420877), (37131,-0.431039), (37132,-0.581943), (37133,-0.622297), (37134,-0.806180), (37135,-0.561799), (37136,-0.725709), (37137,-0.770709), (37138,-0.496600), (37139,-0.347905), (37140,-0.501131), (37141,-0.555420), (37142,-0.613425), (37143,-0.329563), (37144,-0.494401), (37145,-0.637873), (37146,-0.609482), (37147,-0.350702), (37148,-0.432396), (37149,-0.613492), (37150,-0.324520), (37151,-0.488430), (37152,-0.534357), (37153,-0.690371), (37154,-0.569081), (37155,-0.316339), (37156,-0.357158), (37157,-0.520139), (37158,-0.228380), (37159,-0.286385), (37160,-0.624015), (37161,-0.750301), (37162,-0.336844), (37163,-0.486355), (37164,-0.571300), (37165,-0.705947), (37166,-0.466676), (37167,-0.632443), (37168,-0.670011), (37169,-0.787471), (37170,-0.255568), (37171,-0.404150), (37172,-0.489560), (37173,-0.666475), (37174,-0.312009), (37175,-0.477312), (37176,-0.594308), (37177,-0.737780), (37178,-0.354051), (37179,-0.494271), (37180,-0.533232), (37181,-0.719438), (37182,-0.439755), (37183,-0.586478), (37184,-0.633800), (37185,-0.786098), (37186,-0.199384), (37187,-0.379552), (37188,-0.432911), (37189,-0.596357), (37190,-0.228420), (37191,-0.379324), (37192,-0.520009), (37193,-0.669055), (37194,-0.284397), (37195,-0.442733), (37196,-0.518853), (37197,-0.644674), (37198,-0.402151), (37199,-0.553984), (37200,-0.614776), (37201,-0.776828), (37202,-0.226809), (37203,-0.379571), (37204,-0.468698), (37205,-0.627963), (37206,-0.256775), (37207,-0.404892), (37208,-0.415983), (37209,-0.565029), (37210,-0.553359), (37211,-0.310837), (37212,-0.332147), (37213,-0.522997), (37214,-0.225664), (37215,-0.449029), (37216,-0.493563), (37217,-0.629604), (37218,-0.494843), (37219,-0.250927), (37220,-0.299642), (37221,-0.496995), (37222,-0.230319), (37223,-0.298078), (37224,-0.567428), (37225,-0.698359), (37226,-0.310449), (37227,-0.465534), (37228,-0.533293), (37229,-0.673049), (37230,-0.399869), (37231,-0.551703), (37232,-0.611565), (37233,-0.765256), (37234,-0.238462), (37235,-0.332698), (37236,-0.394419), (37237,-0.568548), (37238,-0.251705), (37239,-0.398894), (37240,-0.603214), (37241,-0.735074), (37242,-0.338339), (37243,-0.491566), (37244,-0.553286), (37245,-0.693042), (37246,-0.466312), (37247,-0.601424), (37248,-0.861019), (37249,-0.898122), (37250,-0.652347), (37251,-0.518052), (37252,-0.637370), (37253,-0.721387), (37254,-0.777534), (37255,-0.495064), (37256,-0.674303), (37257,-0.721160), (37258,-0.491643), (37259,-0.439562), (37260,-0.593253), (37261,-0.659619), (37262,-0.824922), (37263,-0.532234), (37264,-0.692428), (37265,-0.763903), (37266,-0.499549), (37267,-0.369434), (37268,-0.552852), (37269,-0.628044), (37270,-0.663753), (37271,-0.398470), (37272,-0.642737), (37273,-0.779706), (37274,-0.434530), (37275,-0.597511), (37276,-0.607673), (37277,-0.719559), (37278,-0.798467), (37279,-0.947513), (37280,-0.670617), (37281,-0.827560), (37282,-0.474487), (37283,-0.643042), (37284,-0.537080), (37285,-0.666153), (37286,-0.612679), (37287,-0.781234), (37288,-0.514557), (37289,-0.669641), (37290,-0.334684), (37291,-0.479549), (37292,-0.500395), (37293,-0.642938), (37294,-0.741819), (37295,-0.877859), (37296,-0.609789), (37297,-0.734681), (37298,-0.409013), (37299,-0.553879), (37300,-0.461852), (37301,-0.580242), (37302,-0.569966), (37303,-0.731553), (37304,-0.699446), (37305,-0.846169), (37306,-0.497742), (37307,-0.617989), (37308,-0.612359), (37309,-0.747469), (37310,-0.828699), (37311,-0.995396), (37312,-0.704101), (37313,-0.842928), (37314,-0.493572), (37315,-0.654694), (37316,-0.524579), (37317,-0.678734), (37318,-0.656382), (37319,-0.799390), (37320,-0.494160), (37321,-0.637632), (37322,-0.289204), (37323,-0.455436), (37324,-0.427510), (37325,-0.597458), (37326,-0.693551), (37327,-0.868145), (37328,-0.571276), (37329,-0.750978), (37330,-0.382113), (37331,-0.514437), (37332,-0.381071), (37333,-0.548696), (37334,-0.507764), (37335,-0.673996), (37336,-0.627490), (37337,-0.763066), (37338,-0.447617), (37339,-0.584586), (37340,-0.582671), (37341,-0.728466), (37342,-0.812947), (37343,-0.926692), (37344,-0.635396), (37345,-0.806738), (37346,-0.435550), (37347,-0.571590), (37348,-0.457732), (37349,-0.603063), (37350,-0.576530), (37351,-0.721395), (37352,-0.470976), (37353,-0.606551), (37354,-0.277168), (37355,-0.431788), (37356,-0.426157), (37357,-0.612362), (37358,-0.643427), (37359,-0.800834), (37360,-0.541125), (37361,-0.699460), (37362,-0.388192), (37363,-0.511226), (37364,-0.389472), (37365,-0.547344), (37366,-0.515236), (37367,-0.645702), (37368,-0.271263), (37369,-0.432850), (37370,-0.451838), (37371,-0.245545), (37372,-0.233876), (37373,-0.384316), (37374,-0.433031), (37375,-0.626204), (37376,-0.327013), (37377,-0.492781), (37378,-0.528490), (37379,-0.292934), (37380,-0.145633), (37381,-0.339734), (37382,-0.375444), (37383,-0.430662), (37384,-0.360002), (37385,-0.517874), (37386,-0.541506), (37387,-0.314311), (37388,-0.299391), (37389,-0.443791), (37390,-0.509693), (37391,-0.746064), (37392,-0.462201), (37393,-0.618214), (37394,-0.658568), (37395,-0.384924), (37396,-0.217185), (37397,-0.359264), (37398,-0.434455), (37399,-0.531942), (37400,-0.473823), (37401,-0.512784), (37402,-0.671120), (37403,-0.235832), (37404,-0.398813), (37405,-0.434987), (37406,-0.605863), (37407,-0.351264), (37408,-0.508671), (37409,-0.566211), (37410,-0.726869), (37411,-0.149446), (37412,-0.299421), (37413,-0.362071), (37414,-0.510188), (37415,-0.138071), (37416,-0.579284), (37417,-0.623354), (37418,-0.395695), (37419,-0.369162), (37420,-0.543755), (37421,-0.580858), (37422,-0.743839), (37423,-0.476233), (37424,-0.651291), (37425,-0.718586), (37426,-0.469560), (37427,-0.310646), (37428,-0.490813), (37429,-0.534419), (37430,-0.569199), (37431,-0.307167), (37432,-0.421840), (37433,-0.432003), (37434,-0.569437), (37435,-0.177810), (37436,-0.323605), (37437,-0.385791), (37438,-0.510218), (37439,-0.292778), (37440,-0.433928), (37441,-0.493791), (37442,-0.680925), (37443,-0.108611), (37444,-0.270663), (37445,-0.350499), (37446,-0.522305), (37447,-0.159014), (37448,-0.419074), (37449,-0.467324), (37450,-0.630305), (37451,-0.220564), (37452,-0.356140), (37453,-0.431796), (37454,-0.540895), (37455,-0.297443), (37456,-0.452992), (37457,-0.505423), (37458,-0.661901), (37459,-0.104915), (37460,-0.288334), (37461,-0.333333), (37462,-0.470302), (37463,-0.079141), (37464,-0.328518), (37465,-0.412535), (37466,-0.547645), (37467,-0.140227), (37468,-0.304602), (37469,-0.394656), (37470,-0.553921), (37471,-0.310005), (37472,-0.484133), (37473,-0.503585), (37474,-0.679572), (37475,-0.089607), (37476,-0.255840), (37477,-0.318954), (37478,-0.465213), (37479,-0.099135), (37480,-0.496685), (37481,-0.546794), (37482,-0.311703), (37483,-0.289815), (37484,-0.417030), (37485,-0.505691), (37486,-0.631512), (37487,-0.383880), (37488,-0.496231), (37489,-0.576067), (37490,-0.339583), (37491,-0.171843), (37492,-0.317638), (37493,-0.381217), (37494,-0.449905), (37495,-0.185086), (37496,-0.602610), (37497,-0.656899), (37498,-0.393010), (37499,-0.381340), (37500,-0.545250), (37501,-0.559593), (37502,-0.736508), (37503,-0.478657), (37504,-0.786560), (37505,-0.841314), (37506,-0.588572), (37507,-0.452883), (37508,-0.624689), (37509,-0.698022), (37510,-0.781110), (37511,-0.450333), (37512,-0.730831), (37513,-0.778153), (37514,-0.513334), (37515,-0.477976), (37516,-0.637240), (37517,-0.727296), (37518,-0.889812), (37519,-0.611523), (37520,-0.794013), (37521,-0.820896), (37522,-0.615068), (37523,-0.477985), (37524,-0.614025), (37525,-0.666921), (37526,-0.709598), (37527,-0.454998), (37528,-0.472127), (37529,-0.646721), (37530,-0.697758), (37531,-0.457094), (37532,-0.458895), (37533,-0.584716), (37534,-0.652011), (37535,-0.851687), (37536,-0.550637), (37537,-0.740095), (37538,-0.777197), (37539,-0.537461), (37540,-0.379941), (37541,-0.551282), (37542,-0.542865), (37543,-0.628275), (37544,-0.565976), (37545,-0.718738), (37546,-0.387497), (37547,-0.512388), (37548,-0.501184), (37549,-0.656268), (37550,-0.739356), (37551,-0.909769), (37552,-0.582244), (37553,-0.732683), (37554,-0.394009), (37555,-0.570925), (37556,-0.428269), (37557,-0.556877), (37558,-0.514087), (37559,-0.672423), (37560,-0.656573), (37561,-0.777749), (37562,-0.447436), (37563,-0.621565), (37564,-0.608038), (37565,-0.799353), (37566,-0.883834), (37567,-1.017087), (37568,-0.719289), (37569,-0.871123), (37570,-0.520837), (37571,-0.676850), (37572,-0.536980), (37573,-0.704142), (37574,-0.657171), (37575,-0.793211), (37576,-0.540469), (37577,-0.677903), (37578,-0.356416), (37579,-0.556557), (37580,-0.552319), (37581,-0.686036), (37582,-0.760299), (37583,-0.910738), (37584,-0.640810), (37585,-0.784747), (37586,-0.441428), (37587,-0.601622), (37588,-0.469649), (37589,-0.594077), (37590,-0.605168), (37591,-0.725880), (37592,-0.433656), (37593,-0.617539), (37594,-0.648603), (37595,-0.435808), (37596,-0.433893), (37597,-0.572256), (37598,-0.643267), (37599,-0.857342), (37600,-0.566047), (37601,-0.724848), (37602,-0.782387), (37603,-0.540794), (37604,-0.349830), (37605,-0.506308), (37606,-0.552700), (37607,-0.621388), (37608,-0.345886), (37609,-0.507474), (37610,-0.594742), (37611,-0.339213), (37612,-0.303855), (37613,-0.452437), (37614,-0.513693), (37615,-0.675280), (37616,-0.439260), (37617,-0.603634), (37618,-0.639808), (37619,-0.392176), (37620,-0.216540), (37621,-0.391597), (37622,-0.433346), (37623,-0.527581), (37624,-0.338939), (37625,-0.474979), (37626,-0.517656), (37627,-0.284888), (37628,-0.263464), (37629,-0.421800), (37630,-0.480734), (37631,-0.642786), (37632,-0.414198), (37633,-0.558134), (37634,-0.597559), (37635,-0.349463), (37636,-0.214238), (37637,-0.384186), (37638,-0.391561), (37639,-0.472791), (37640,-0.357539), (37641,-0.529345), (37642,-0.610111), (37643,-0.324390), (37644,-0.323869), (37645,-0.471057), (37646,-0.555538), (37647,-0.758930), (37648,-0.464848), (37649,-0.612500), (37650,-0.649603), (37651,-0.403829), (37652,-0.246308), (37653,-0.405573), (37654,-0.431064), (37655,-0.464915), (37656,-0.548467), (37657,-0.596253), (37658,-0.746692), (37659,-0.336952), (37660,-0.486927), (37661,-0.558402), (37662,-0.736711), (37663,-0.496046), (37664,-0.649737), (37665,-0.698917), (37666,-0.846569), (37667,-0.280758), (37668,-0.429339), (37669,-0.485951), (37670,-0.663796), (37671,-0.283318), (37672,-0.425397), (37673,-0.498265), (37674,-0.616190), (37675,-0.216203), (37676,-0.396835), (37677,-0.490141), (37678,-0.650335), (37679,-0.410135), (37680,-0.522486), (37681,-0.594890), (37682,-0.736040), (37683,-0.178589), (37684,-0.350860), (37685,-0.387499), (37686,-0.560233), (37687,-0.184865), (37688,-0.444925), (37689,-0.490854), (37690,-0.643151), (37691,-0.239913), (37692,-0.395927), (37693,-0.460899), (37694,-0.606693), (37695,-0.366028), (37696,-0.479308), (37697,-0.549390), (37698,-0.703081), (37699,-0.175823), (37700,-0.308611), (37701,-0.394486), (37702,-0.530062), (37703,-0.169093), (37704,-0.431011), (37705,-0.535465), (37706,-0.697517), (37707,-0.282667), (37708,-0.430784), (37709,-0.512942), (37710,-0.646196), (37711,-0.380912), (37712,-0.529958), (37713,-0.559165), (37714,-0.716107), (37715,-0.142864), (37716,-0.296091), (37717,-0.377784), (37718,-0.497567), (37719,-0.155643), (37720,-0.508137), (37721,-0.594012), (37722,-0.771392), (37723,-0.373728), (37724,-0.507910), (37725,-0.553838), (37726,-0.678266), (37727,-0.444104), (37728,-0.620090), (37729,-0.711539), (37730,-0.829928), (37731,-0.290594), (37732,-0.467974), (37733,-0.543630), (37734,-0.721474), (37735,-0.362827), (37736,-0.603379), (37737,-0.636766), (37738,-0.395636), (37739,-0.370497), (37740,-0.530691), (37741,-0.578012), (37742,-0.729381), (37743,-0.490573), (37744,-0.608034), (37745,-0.659536), (37746,-0.430948), (37747,-0.278073), (37748,-0.447092), (37749,-0.464221), (37750,-0.564495), (37751,-0.216996), (37752,-0.621050), (37753,-0.689274), (37754,-0.459757), (37755,-0.463881), (37756,-0.601314), (37757,-0.703910), (37758,-0.900800), (37759,-0.600214), (37760,-0.708850), (37761,-0.751991), (37762,-0.910327), (37763,-0.371920), (37764,-0.540475), (37765,-0.583617), (37766,-0.730340), (37767,-0.414891), (37768,-0.538855), (37769,-0.704158), (37770,-0.757054), (37771,-0.488519), (37772,-0.421575), (37773,-0.626825), (37774,-0.629090), (37775,-0.834340), (37776,-0.566734), (37777,-0.720890), (37778,-0.776108), (37779,-0.547520), (37780,-0.374206), (37781,-0.510247), (37782,-0.558497), (37783,-0.657378), (37784,-0.504038), (37785,-0.636826), (37786,-0.671607), (37787,-0.445806), (37788,-0.460613), (37789,-0.585969), (37790,-0.626788), (37791,-0.809742), (37792,-0.528202), (37793,-0.682821), (37794,-0.768232), (37795,-0.512703), (37796,-0.357040), (37797,-0.505622), (37798,-0.582207), (37799,-0.677371), (37800,-0.637368), (37801,-0.767834), (37802,-0.450528), (37803,-0.580065), (37804,-0.565609), (37805,-0.712797), (37806,-0.779163), (37807,-0.910558), (37808,-0.634127), (37809,-0.782244), (37810,-0.472834), (37811,-0.592152), (37812,-0.466681), (37813,-0.644526), (37814,-0.603594), (37815,-0.728486), (37816,-0.492466), (37817,-0.663808), (37818,-0.741322), (37819,-0.502515), (37820,-0.489916), (37821,-0.665439), (37822,-0.682568), (37823,-0.845084), (37824,-0.571905), (37825,-0.777619), (37826,-0.790568), (37827,-0.567554), (37828,-0.421646), (37829,-0.601349), (37830,-0.624516), (37831,-0.715036), (37832,-0.459507), (37833,-0.628526), (37834,-0.674919), (37835,-0.421713), (37836,-0.379387), (37837,-0.543761), (37838,-0.613379), (37839,-0.803765), (37840,-0.509219), (37841,-0.662909), (37842,-0.715340), (37843,-0.436122), (37844,-0.299969), (37845,-0.436474), (37846,-0.487975), (37847,-0.585462), (37848,-0.464173), (37849,-0.654558), (37850,-0.719531), (37851,-0.475150), (37852,-0.456978), (37853,-0.646435), (37854,-0.701653), (37855,-0.869743), (37856,-0.578913), (37857,-0.733068), (37858,-0.808259), (37859,-0.602896), (37860,-0.421222), (37861,-0.570732), (37862,-0.588327), (37863,-0.677917), (37864,-0.393590), (37865,-0.550068), (37866,-0.589493), (37867,-0.320958), (37868,-0.315792), (37869,-0.477844), (37870,-0.534455), (37871,-0.691397), (37872,-0.409393), (37873,-0.551471), (37874,-0.630378), (37875,-0.365095), (37876,-0.255418), (37877,-0.418863), (37878,-0.472223), (37879,-0.536731), (37880,-0.417299), (37881,-0.567739), (37882,-0.633640), (37883,-0.382756), (37884,-0.369694), (37885,-0.496444), (37886,-0.538191), (37887,-0.765272), (37888,-0.465617), (37889,-0.632314), (37890,-0.683816), (37891,-0.436648), (37892,-0.245684), (37893,-0.423064), (37894,-0.473637), (37895,-0.525604), (37896,-0.409888), (37897,-0.562185), (37898,-0.616474), (37899,-0.418542), (37900,-0.413841), (37901,-0.602369), (37902,-0.647832), (37903,-0.820568), (37904,-0.500474), (37905,-0.677854), (37906,-0.741433), (37907,-0.508665), (37908,-0.372511), (37909,-0.516912), (37910,-0.580026), (37911,-0.616200), (37912,-0.411766), (37913,-0.435863), (37914,-0.603489), (37915,-0.580207), (37916,-0.324213), (37917,-0.383148), (37918,-0.556347), (37919,-0.291064), (37920,-0.502353), (37921,-0.557571), (37922,-0.691752), (37923,-0.546774), (37924,-0.287064), (37925,-0.385016), (37926,-0.546139), (37927,-0.228368), (37928,-0.505614), (37929,-0.588702), (37930,-0.673647), (37931,-0.282022), (37932,-0.425494), (37933,-0.476532), (37934,-0.657163), (37935,-0.407208), (37936,-0.529778), (37937,-0.582673), (37938,-0.717784), (37939,-0.168231), (37940,-0.321922), (37941,-0.386894), (37942,-0.518289), (37943,-0.183796), (37944,-0.519569), (37945,-0.596618), (37946,-0.739162), (37947,-0.350323), (37948,-0.511910), (37949,-0.551800), (37950,-0.717103), (37951,-0.454607), (37952,-0.603653), (37953,-0.644007), (37954,-0.792588), (37955,-0.212378), (37956,-0.357708), (37957,-0.484922), (37958,-0.627466), (37959,-0.236304), (37960,-0.481501), (37961,-0.550189), (37962,-0.710383), (37963,-0.306216), (37964,-0.460836), (37965,-0.542066), (37966,-0.688325), (37967,-0.434654), (37968,-0.569300), (37969,-0.633344), (37970,-0.781925), (37971,-0.250022), (37972,-0.398139), (37973,-0.445461), (37974,-0.574069), (37975,-0.232609), (37976,-0.316625), (37977,-0.405752), (37978,-0.586383), (37979,-0.576572), (37980,-0.323366), (37981,-0.388338), (37982,-0.512766), (37983,-0.225187), (37984,-0.443908), (37985,-0.488442), (37986,-0.650494), (37987,-0.489722), (37988,-0.267172), (37989,-0.307062), (37990,-0.450534), (37991,-0.139266), (37992,-0.423479), (37993,-0.587854), (37994,-0.242678), (37995,-0.387078), (37996,-0.388415), (37997,-0.530030), (37998,-0.642381), (37999,-0.773311), (38000,-0.484803), (38001,-0.627346), (38002,-0.298892), (38003,-0.428429), (38004,-0.291811), (38005,-0.451540), (38006,-0.436619), (38007,-0.609355), (38008,-0.467627), (38009,-0.497297), (38010,-0.668175), (38011,-0.251467), (38012,-0.394939), (38013,-0.449692), (38014,-0.591306), (38015,-0.352963), (38016,-0.521519), (38017,-0.692395), (38018,-0.720673), (38019,-0.491620), (38020,-0.346642), (38021,-0.509622), (38022,-0.566234), (38023,-0.604730), (38024,-0.479724), (38025,-0.614835), (38026,-0.654261), (38027,-0.403841), (38028,-0.380560), (38029,-0.570945), (38030,-0.635918), (38031,-0.808653), (38032,-0.530364), (38033,-0.697525), (38034,-0.752279), (38035,-0.534839), (38036,-0.357345), (38037,-0.535190), (38038,-0.600162), (38039,-0.659096), (38040,-0.583326), (38041,-0.748165), (38042,-0.769011), (38043,-0.550642), (38044,-0.504135), (38045,-0.647143), (38046,-0.716296), (38047,-0.925726), (38048,-0.640005), (38049,-0.792302), (38050,-0.815470), (38051,-0.589205), (38052,-0.444225), (38053,-0.570047), (38054,-0.616439), (38055,-0.684664), (38056,-0.766358), (38057,-0.503397), (38058,-0.659875), (38059,-0.331420), (38060,-0.503691), (38061,-0.497132), (38062,-0.680085), (38063,-0.738091), (38064,-0.896891), (38065,-0.583300), (38066,-0.708192), (38067,-0.328179), (38068,-0.505559), (38069,-0.349897), (38070,-0.496155), (38071,-0.475197), (38072,-0.500687), (38073,-0.634404), (38074,-0.688229), (38075,-0.435952), (38076,-0.436360), (38077,-0.596553), (38078,-0.646662), (38079,-0.843551), (38080,-0.572694), (38081,-0.700373), (38082,-0.759307), (38083,-0.506565), (38084,-0.382953), (38085,-0.534321), (38086,-0.613693), (38087,-0.673556), (38088,-0.756180), (38089,-0.476961), (38090,-0.632510), (38091,-0.288728), (38092,-0.412226), (38093,-0.414957), (38094,-0.578866), (38095,-0.646626), (38096,-0.773376), (38097,-0.504841), (38098,-0.683150), (38099,-0.337045), (38100,-0.481910), (38101,-0.363872), (38102,-0.469720), (38103,-0.484063), (38104,-0.557396), (38105,-0.693436), (38106,-0.762589), (38107,-0.538181), (38108,-0.539054), (38109,-0.673236), (38110,-0.739137), (38111,-0.881216), (38112,-0.637299), (38113,-0.787274), (38114,-0.867575), (38115,-0.639451), (38116,-0.493078), (38117,-0.665814), (38118,-0.718245), (38119,-0.730265), (38120,-0.810566), (38121,-0.537850), (38122,-0.651595), (38123,-0.331966), (38124,-0.475903), (38125,-0.476775), (38126,-0.643936), (38127,-0.722379), (38128,-0.879321), (38129,-0.580130), (38130,-0.729641), (38131,-0.411869), (38132,-0.560451), (38133,-0.430335), (38134,-0.585420), (38135,-0.522192), (38136,-0.424591), (38137,-0.554593), (38138,-0.620958), (38139,-0.359392), (38140,-0.361657), (38141,-0.482369), (38142,-0.543161), (38143,-0.738656), (38144,-0.479876), (38145,-0.631709), (38146,-0.701791), (38147,-0.460662), (38148,-0.312431), (38149,-0.477270), (38150,-0.518089), (38151,-0.622543), (38152,-0.818038), (38153,-0.548110), (38154,-0.666035), (38155,-0.325039), (38156,-0.443893), (38157,-0.440584), (38158,-0.594740), (38159,-0.692692), (38160,-0.848705), (38161,-0.556946), (38162,-0.707385), (38163,-0.373821), (38164,-0.541447), (38165,-0.406222), (38166,-0.544121), (38167,-0.521768), (38168,-0.290392), (38169,-0.423182), (38170,-0.493264), (38171,-0.686901), (38172,-0.258580), (38173,-0.374182), (38174,-0.453554), (38175,-0.615141), (38176,-0.390269), (38177,-0.514232), (38178,-0.585244), (38179,-0.758908), (38180,-0.220502), (38181,-0.357006), (38182,-0.406186), (38183,-0.553838), (38184,-0.461347), (38185,-0.568589), (38186,-0.660966), (38187,-0.458390), (38188,-0.443469), (38189,-0.600876), (38190,-0.628225), (38191,-0.797708), (38192,-0.497123), (38193,-0.655924), (38194,-0.744121), (38195,-0.502992), (38196,-0.351045), (38197,-0.509381), (38198,-0.542303), (38199,-0.597057), (38200,-0.423743), (38201,-0.608091), (38202,-0.677244), (38203,-0.424037), (38204,-0.423051), (38205,-0.570240), (38206,-0.619884), (38207,-0.826991), (38208,-0.534767), (38209,-0.702858), (38210,-0.727884), (38211,-0.469568), (38212,-0.306009), (38213,-0.463416), (38214,-0.500055), (38215,-0.585929), (38216,-0.403791), (38217,-0.558410), (38218,-0.621989), (38219,-0.383182), (38220,-0.337605), (38221,-0.495941), (38222,-0.549765), (38223,-0.728075), (38224,-0.454430), (38225,-0.628094), (38226,-0.684242), (38227,-0.448221), (38228,-0.277695), (38229,-0.395620), (38230,-0.476385), (38231,-0.514882), (38232,-0.218942), (38233,-0.380529), (38234,-0.456649), (38235,-0.640997), (38236,-0.240546), (38237,-0.366367), (38238,-0.429017), (38239,-0.535330), (38240,-0.304883), (38241,-0.432098), (38242,-0.503573), (38243,-0.661909), (38244,-0.117000), (38245,-0.268369), (38246,-0.337986), (38247,-0.486103), (38248,-0.396399), (38249,-0.531975), (38250,-0.588122), (38251,-0.345598), (38252,-0.342291), (38253,-0.490408), (38254,-0.503821), (38255,-0.708142), (38256,-0.405234), (38257,-0.565428), (38258,-0.607640), (38259,-0.346538), (38260,-0.184837), (38261,-0.360823), (38262,-0.403965), (38263,-0.464757), (38264,-0.345325), (38265,-0.534318), (38266,-0.612296), (38267,-0.415293), (38268,-0.391083), (38269,-0.517368), (38270,-0.551684), (38271,-0.725813), (38272,-0.484684), (38273,-0.672282), (38274,-0.716817), (38275,-0.490551), (38276,-0.331637), (38277,-0.474645), (38278,-0.512212), (38279,-0.595300), (38280,-0.447999), (38281,-0.610515), (38282,-0.629966), (38283,-0.394876), (38284,-0.351621), (38285,-0.514137), (38286,-0.591651), (38287,-0.782037), (38288,-0.467053), (38289,-0.663013), (38290,-0.716373), (38291,-0.448767), (38292,-0.295892), (38293,-0.474665), (38294,-0.495975), (38295,-0.582779), (38296,-0.832156), (38297,-0.555260), (38298,-0.750756), (38299,-0.419050), (38300,-0.532330), (38301,-0.537846), (38302,-0.664597), (38303,-0.741182), (38304,-0.899982), (38305,-0.591036), (38306,-0.720109), (38307,-0.391190), (38308,-0.536056), (38309,-0.401295), (38310,-0.561025), (38311,-0.556323), (38312,-0.911604), (38313,-0.610091), (38314,-0.361994), (38315,-0.423715), (38316,-0.582051), (38317,-0.569453), (38318,-0.733363), (38319,-0.767678), (38320,-0.898145), (38321,-0.617533), (38322,-0.386158), (38323,-0.426048), (38324,-0.602034), (38325,-0.492357), (38326,-0.566619), (38327,-0.607438), (38328,-0.787140), (38329,-0.504207), (38330,-0.671368), (38331,-0.316902), (38332,-0.459444), (38333,-0.509553), (38334,-0.673463), (38335,-0.728216), (38336,-0.830349), (38337,-0.559956), (38338,-0.708073), (38339,-0.357787), (38340,-0.544922), (38341,-0.391117), (38342,-0.535054), (38343,-0.507127), (38344,-0.705409), (38345,-0.419224), (38346,-0.547368), (38347,-0.207301), (38348,-0.383288), (38349,-0.342356), (38350,-0.504407), (38351,-0.588889), (38352,-0.734683), (38353,-0.426201), (38354,-0.580822), (38355,-0.249580), (38356,-0.367041), (38357,-0.261079), (38358,-0.430563), (38359,-0.397062), (38360,-0.782536), (38361,-0.553948), (38362,-0.697420), (38363,-0.372681), (38364,-0.533340), (38365,-0.493801), (38366,-0.643776), (38367,-0.728257), (38368,-0.875445), (38369,-0.625490), (38370,-0.778717), (38371,-0.421928), (38372,-0.557968), (38373,-0.408808), (38374,-0.595943), (38375,-0.546649), (38376,-0.705915), (38377,-0.432735), (38378,-0.582245), (38379,-0.256114), (38380,-0.413985), (38381,-0.441798), (38382,-0.573193), (38383,-0.641881), (38384,-0.780244), (38385,-0.520999), (38386,-0.662148), (38387,-0.303967), (38388,-0.475308), (38389,-0.312678), (38390,-0.480769), (38391,-0.466313), (38392,-0.656234), (38393,-0.386306), (38394,-0.520488), (38395,-0.186924), (38396,-0.339686), (38397,-0.360996), (38398,-0.483101), (38399,-0.541106), (38400,-0.679469), (38401,-0.437410), (38402,-0.569270), (38403,-0.268686), (38404,-0.403332), (38405,-0.271358), (38406,-0.413437), (38407,-0.346958), (38408,-0.696201), (38409,-0.413732), (38410,-0.587396), (38411,-0.210633), (38412,-0.401948), (38413,-0.387028), (38414,-0.526319), (38415,-0.579680), (38416,-0.773782), (38417,-0.470874), (38418,-0.607379), (38419,-0.289608), (38420,-0.419145), (38421,-0.291817), (38422,-0.440862), (38423,-0.402717), (38424,-0.195032), (38425,-0.322710), (38426,-0.416946), (38427,-0.559954), (38428,-0.148819), (38429,-0.274640), (38430,-0.313137), (38431,-0.458003), (38432,-0.218731), (38433,-0.372886), (38434,-0.430427), (38435,-0.597123), (38436,-0.054537), (38437,-0.204047), (38438,-0.272272), (38439,-0.399486), (38440,-0.284699), (38441,-0.423991), (38442,-0.495931), (38443,-0.249227), (38444,-0.269144), (38445,-0.405184), (38446,-0.449254), (38447,-0.606196), (38448,-0.337662), (38449,-0.524796), (38450,-0.608348), (38451,-0.354677), (38452,-0.208305), (38453,-0.381969), (38454,-0.419072), (38455,-0.499837), (38456,-0.307015), (38457,-0.462100), (38458,-0.514531), (38459,-0.277117), (38460,-0.307252), (38461,-0.436790), (38462,-0.472034), (38463,-0.643376), (38464,-0.375771), (38465,-0.540145), (38466,-0.565171), (38467,-0.348195), (38468,-0.192068), (38469,-0.385705), (38470,-0.435349), (38471,-0.498464), (38472,-0.309822), (38473,-0.437502), (38474,-0.488075), (38475,-0.261809), (38476,-0.263146), (38477,-0.438668), (38478,-0.492493), (38479,-0.681485), (38480,-0.378113), (38481,-0.490464), (38482,-0.554043), (38483,-0.317558), (38484,-0.215313), (38485,-0.392693), (38486,-0.454414), (38487,-0.524032), (38488,-0.154701), (38489,-0.310715), (38490,-0.352927), (38491,-0.524269), (38492,-0.130321), (38493,-0.256606), (38494,-0.321579), (38495,-0.438575), (38496,-0.180724), (38497,-0.359497), (38498,-0.428650), (38499,-0.576767), (38500,-0.035574), (38501,-0.191123), (38502,-0.249593), (38503,-0.412573), (38504,-0.416697), (38505,-0.566207), (38506,-0.236824), (38507,-0.390050), (38508,-0.357479), (38509,-0.510241), (38510,-0.582181), (38511,-0.738658), (38512,-0.485917), (38513,-0.614525), (38514,-0.279103), (38515,-0.424433), (38516,-0.296176), (38517,-0.406669), (38518,-0.398251), (38519,-0.524072), (38520,-0.242996), (38521,-0.402725), (38522,-0.475595), (38523,-0.225639), (38524,-0.220938), (38525,-0.404356), (38526,-0.489766), (38527,-0.628129), (38528,-0.514271), (38529,-0.644737), (38530,-0.722716), (38531,-0.480657), (38532,-0.330104), (38533,-0.500053), (38534,-0.555270), (38535,-0.613740), (38536,-0.434853), (38537,-0.580647), (38538,-0.596383), (38539,-0.378014), (38540,-0.364487), (38541,-0.502849), (38542,-0.556209), (38543,-0.753098), (38544,-0.463197), (38545,-0.600166), (38546,-0.656778), (38547,-0.427260), (38548,-0.271598), (38549,-0.427612), (38550,-0.487010), (38551,-0.598432), (38552,-0.847809), (38553,-0.565804), (38554,-0.752474), (38555,-0.377105), (38556,-0.575387), (38557,-0.567435), (38558,-0.696972), (38559,-0.764731), (38560,-0.909132), (38561,-0.591361), (38562,-0.732975), (38563,-0.386870), (38564,-0.507581), (38565,-0.385363), (38566,-0.560885), (38567,-0.518559), (38568,-0.708945), (38569,-0.465493), (38570,-0.607107), (38571,-0.295374), (38572,-0.440240), (38573,-0.436467), (38574,-0.605951), (38575,-0.691825), (38576,-0.851555), (38577,-0.569086), (38578,-0.692120), (38579,-0.388748), (38580,-0.518285), (38581,-0.390028), (38582,-0.545112), (38583,-0.480955), (38584,-0.831592), (38585,-0.572347), (38586,-0.720928), (38587,-0.349741), (38588,-0.482065), (38589,-0.525671), (38590,-0.650563), (38591,-0.745727), (38592,-0.919391), (38593,-0.664327), (38594,-0.804548), (38595,-0.448688), (38596,-0.572187), (38597,-0.428601), (38598,-0.544668), (38599,-0.529283), (38600,-0.731746), (38601,-0.464140), (38602,-0.624334), (38603,-0.293093), (38604,-0.447248), (38605,-0.443940), (38606,-0.588340), (38607,-0.669570), (38608,-0.820010), (38609,-0.534754), (38610,-0.680084), (38611,-0.346984), (38612,-0.513681), (38613,-0.386352), (38614,-0.507993), (38615,-0.465667), (38616,-0.855786), (38617,-0.594683), (38618,-0.754413), (38619,-0.410165), (38620,-0.586617), (38621,-0.582844), (38622,-0.704020), (38623,-0.785715), (38624,-0.950553), (38625,-0.679231), (38626,-0.825026), (38627,-0.487282), (38628,-0.594523), (38629,-0.466731), (38630,-0.613454), (38631,-0.623151), (38632,-0.786597), (38633,-0.489263), (38634,-0.635523), (38635,-0.317287), (38636,-0.452398), (38637,-0.455593), (38638,-0.598136), (38639,-0.698410), (38640,-0.866035), (38641,-0.589604), (38642,-0.720535), (38643,-0.363282), (38644,-0.510934), (38645,-0.376174), (38646,-0.556806), (38647,-0.540027), (38648,-0.683963), (38649,-0.434938), (38650,-0.572836), (38651,-0.247169), (38652,-0.372990), (38653,-0.391512), (38654,-0.517334), (38655,-0.605067), (38656,-0.704411), (38657,-0.400111), (38658,-0.539402), (38659,-0.214664), (38660,-0.394831), (38661,-0.251245), (38662,-0.394717), (38663,-0.393732), (38664,-0.705815), (38665,-0.420095), (38666,-0.554741), (38667,-0.217926), (38668,-0.414815), (38669,-0.371095), (38670,-0.509923), (38671,-0.581862), (38672,-0.728586), (38673,-0.433111), (38674,-0.594233), (38675,-0.255095), (38676,-0.452449), (38677,-0.293999), (38678,-0.436542), (38679,-0.439273), (38680,-0.195820), (38681,-0.350905), (38682,-0.438173), (38683,-0.567711), (38684,-0.167259), (38685,-0.342317), (38686,-0.389174), (38687,-0.544258), (38688,-0.273401), (38689,-0.433595), (38690,-0.511574), (38691,-0.647149), (38692,-0.141258), (38693,-0.293555), (38694,-0.355740), (38695,-0.497355), (38696,-0.416011), (38697,-0.570167), (38698,-0.593799), (38699,-0.370785), (38700,-0.367941), (38701,-0.524883), (38702,-0.568489), (38703,-0.728218), (38704,-0.448071), (38705,-0.609195), (38706,-0.676025), (38707,-0.427928), (38708,-0.256473), (38709,-0.372075), (38710,-0.458879), (38711,-0.545682), (38712,-0.348680), (38713,-0.524666), (38714,-0.562234), (38715,-0.350832), (38716,-0.346595), (38717,-0.495640), (38718,-0.519737), (38719,-0.693401), (38720,-0.423938), (38721,-0.596673), (38722,-0.631918), (38723,-0.389395), (38724,-0.229088), (38725,-0.408326), (38726,-0.463079), (38727,-0.542916), (38728,-0.352880), (38729,-0.547447), (38730,-0.559931), (38731,-0.345278), (38732,-0.316887), (38733,-0.513312), (38734,-0.529048), (38735,-0.692493), (38736,-0.416062), (38737,-0.548386), (38738,-0.599423), (38739,-0.363404), (38740,-0.185910), (38741,-0.368864), (38742,-0.450093), (38743,-0.502989), (38744,-0.158277), (38745,-0.358418), (38746,-0.375547), (38747,-0.527381), (38748,-0.102775), (38749,-0.272259), (38750,-0.337232), (38751,-0.483955), (38752,-0.196376), (38753,-0.348209), (38754,-0.418756), (38755,-0.588239), (38756,-0.001526), (38757,-0.151965), (38758,-0.233660), (38759,-0.372487), (38760,-0.194528), (38761,-0.352864), (38762,-0.410869), (38763,-0.152089), (38764,-0.148781), (38765,-0.318265), (38766,-0.360477), (38767,-0.541573), (38768,-0.267464), (38769,-0.428587), (38770,-0.496811), (38771,-0.251965), (38772,-0.098161), (38773,-0.242097), (38774,-0.279665), (38775,-0.385048), (38776,-0.257256), (38777,-0.430920), (38778,-0.516794), (38779,-0.275665), (38780,-0.250061), (38781,-0.387030), (38782,-0.412056), (38783,-0.584326), (38784,-0.553148), (38785,-0.699872), (38786,-0.759735), (38787,-0.507922), (38788,-0.357834), (38789,-0.538001), (38790,-0.583929), (38791,-0.638683), (38792,-0.468156), (38793,-0.640891), (38794,-0.703542), (38795,-0.453122), (38796,-0.464213), (38797,-0.660173), (38798,-0.666619), (38799,-0.834245), (38800,-0.570355), (38801,-0.717543), (38802,-0.774620), (38803,-0.531632), (38804,-0.337416), (38805,-0.511080), (38806,-0.570943), (38807,-0.632665), (38808,-0.772421), (38809,-0.489951), (38810,-0.669189), (38811,-0.315652), (38812,-0.459124), (38813,-0.471144), (38814,-0.600681), (38815,-0.659616), (38816,-0.851394), (38817,-0.613052), (38818,-0.733300), (38819,-0.416922), (38820,-0.592444), (38821,-0.435853), (38822,-0.570964), (38823,-0.523529), (38824,-0.714379), (38825,-0.450489), (38826,-0.566556), (38827,-0.241353), (38828,-0.403405), (38829,-0.403813), (38830,-0.530099), (38831,-0.588568), (38832,-0.708815), (38833,-0.455609), (38834,-0.612551), (38835,-0.286884), (38836,-0.444755), (38837,-0.320678), (38838,-0.458112), (38839,-0.403245), (38840,-0.818446), (38841,-0.532725), (38842,-0.701280), (38843,-0.381651), (38844,-0.541845), (38845,-0.543646), (38846,-0.683866), (38847,-0.749768), (38848,-0.902065), (38849,-0.608448), (38850,-0.756100), (38851,-0.394202), (38852,-0.559041), (38853,-0.424281), (38854,-0.613273), (38855,-0.577450), (38856,-0.725103), (38857,-0.461214), (38858,-0.615833), (38859,-0.261367), (38860,-0.419238), (38861,-0.422897), (38862,-0.574731), (38863,-0.675005), (38864,-0.811509), (38865,-0.529968), (38866,-0.688769), (38867,-0.337555), (38868,-0.523295), (38869,-0.335118), (38870,-0.476268), (38871,-0.461347), (38872,-0.770644), (38873,-0.484458), (38874,-0.668341), (38875,-0.310159), (38876,-0.445735), (38877,-0.429885), (38878,-0.588686), (38879,-0.678741), (38880,-0.818961), (38881,-0.602915), (38882,-0.724555), (38883,-0.396566), (38884,-0.530748), (38885,-0.403884), (38886,-0.582657), (38887,-0.579349), (38888,-0.741865), (38889,-0.469615), (38890,-0.591720), (38891,-0.220532), (38892,-0.389551), (38893,-0.427118), (38894,-0.574307), (38895,-0.642530), (38896,-0.798544), (38897,-0.523042), (38898,-0.670230), (38899,-0.294861), (38900,-0.454126), (38901,-0.326334), (38902,-0.500927), (38903,-0.501334), (38904,-0.511961), (38905,-0.216021), (38906,-0.394795), (38907,-0.463948), (38908,-0.218637), (38909,-0.172132), (38910,-0.316997), (38911,-0.407516), (38912,-0.843156), (38913,-1.001956), (38914,-0.714841), (38915,-0.502975), (38916,-0.555406), (38917,-0.707704), (38918,-0.552041), (38919,-0.635129), (38920,-0.826908), (38921,-0.896990), (38922,-1.036746), (38923,-0.367353), (38924,-0.523831), (38925,-0.596235), (38926,-0.740172), (38927,-0.767056), (38928,-0.892412), (38929,-0.923941), (38930,-1.084600), (38931,-0.435644), (38932,-0.583761), (38933,-0.629689), (38934,-0.785702), (38935,-0.525528), (38936,-0.922150), (38937,-0.668479), (38938,-0.771076), (38939,-0.451911), (38940,-0.587952), (38941,-0.608332), (38942,-0.768061), (38943,-0.853008), (38944,-1.036426), (38945,-0.744202), (38946,-0.877920), (38947,-0.555968), (38948,-0.732883), (38949,-0.563286), (38950,-0.738809), (38951,-0.734572), (38952,-0.785144), (38953,-0.914682), (38954,-0.644754), (38955,-0.375290), (38956,-0.403103), (38957,-0.581876), (38958,-0.589252), (38959,-0.758735), (38960,-0.778651), (38961,-0.907724), (38962,-0.643835), (38963,-0.406886), (38964,-0.479290), (38965,-0.632516), (38966,-0.473138), (38967,-0.567373), (38968,-0.924049), (38969,-0.632754), (38970,-0.797128), (38971,-0.477499), (38972,-0.648376), (38973,-0.604657), (38974,-0.767173), (38975,-0.840971), (38976,-1.006739), (38977,-0.694541), (38978,-0.837549), (38979,-0.495160), (38980,-0.685081), (38981,-0.574011), (38982,-0.673820), (38983,-0.626384), (38984,-0.760103), (38985,-0.911006), (38986,-0.651297), (38987,-0.414813), (38988,-0.468172), (38989,-0.638585), (38990,-0.628774), (38991,-0.828914), (38992,-0.887384), (38993,-1.051294), (38994,-0.768360), (38995,-0.525372), (38996,-0.577804), (38997,-0.724063), (38998,-0.549820), (38999,-0.594820), (39000,-0.907368), (39001,-0.623040), (39002,-0.791130), (39003,-0.461282), (39004,-0.597787), (39005,-0.642786), (39006,-0.763033), (39007,-0.832186), (39008,-0.967297), (39009,-0.695976), (39010,-0.846415), (39011,-0.497059), (39012,-0.674438), (39013,-0.513666), (39014,-0.710091), (39015,-0.667765), (39016,-0.910175), (39017,-1.047608), (39018,-0.392614), (39019,-0.578355), (39020,-0.606168), (39021,-0.759859), (39022,-0.776989), (39023,-0.885623), (39024,-0.973820), (39025,-1.112183), (39026,-0.455796), (39027,-0.655007), (39028,-0.656808), (39029,-0.808641), (39030,-0.562402), (39031,-0.733279), (39032,-0.811258), (39033,-0.940794), (39034,-0.641603), (39035,-0.388862), (39036,-0.470556), (39037,-0.607061), (39038,-0.603288), (39039,-0.758372), (39040,-1.029116), (39041,-1.183271), (39042,-0.496691), (39043,-0.655492), (39044,-0.725574), (39045,-0.894593), (39046,-0.659502), (39047,-0.832237), (39048,-0.997076), (39049,-1.155876), (39050,-0.471155), (39051,-0.596976), (39052,-0.672167), (39053,-0.820284), (39054,-0.829517), (39055,-0.986459), (39056,-1.007769), (39057,-1.159602), (39058,-0.471164), (39059,-0.647615), (39060,-0.713981), (39061,-0.871388), (39062,-0.611215), (39063,-0.806710), (39064,-1.040294), (39065,-1.200488), (39066,-0.530166), (39067,-0.688966), (39068,-0.721888), (39069,-0.876043), (39070,-0.861123), (39071,-1.018065), (39072,-1.082109), (39073,-1.269243), (39074,-0.638403), (39075,-0.779088), (39076,-0.834771), (39077,-0.942012), (39078,-0.719927), (39079,-0.887088), (39080,-0.962279), (39081,-1.003098), (39082,-0.763826), (39083,-0.472532), (39084,-0.628545), (39085,-0.701414), (39086,-0.867181), (39087,-0.830430), (39088,-0.990159), (39089,-1.026333), (39090,-0.807499), (39091,-0.538036), (39092,-0.701945), (39093,-0.733474), (39094,-0.817026), (39095,-0.650216), (39096,-0.973447), (39097,-1.151292), (39098,-0.476789), (39099,-0.625835), (39100,-0.701026), (39101,-0.817558), (39102,-0.842584), (39103,-1.005100), (39104,-1.056602), (39105,-1.181959), (39106,-0.542758), (39107,-0.667185), (39108,-0.757706), (39109,-0.900715), (39110,-0.635431), (39111,-0.798408), (39112,-0.909833), (39113,-0.952042), (39114,-0.705343), (39115,-0.426590), (39116,-0.567739), (39117,-0.649897), (39118,-0.830525), (39119,-0.822108), (39120,-0.985555), (39121,-1.039842), (39122,-0.802429), (39123,-0.517177), (39124,-0.668075), (39125,-0.696821), (39126,-0.765046), (39127,-0.640500), (39128,-1.042698), (39129,-1.216364), (39130,-0.523277), (39131,-0.687187), (39132,-0.744730), (39133,-0.867764), (39134,-0.905332), (39135,-1.049268), (39136,-1.086836), (39137,-1.237741), (39138,-0.586462), (39139,-0.736897), (39140,-0.766106), (39141,-0.917474), (39142,-0.700036), (39143,-0.835612), (39144,-0.914520), (39145,-0.956728), (39146,-0.744400), (39147,-0.445209), (39148,-0.630484), (39149,-0.647614), (39150,-0.845431), (39151,-0.825399), (39152,-0.978163), (39153,-1.029664), (39154,-0.796434), (39155,-0.492597), (39156,-0.654184), (39157,-0.710794), (39158,-0.756258), (39159,-0.614993), (39160,-0.736174), (39161,-0.920985), (39162,-0.288285), (39163,-0.427575), (39164,-0.518098), (39165,-0.667606), (39166,-0.645257), (39167,-0.837964), (39168,-0.909440), (39169,-1.038510), (39170,-0.363080), (39171,-0.497723), (39172,-0.589637), (39173,-0.780954), (39174,-0.498019), (39175,-0.642887), (39176,-0.863929), (39177,-0.947014), (39178,-0.684986), (39179,-0.401124), (39180,-0.565961), (39181,-0.640223), (39182,-0.830144), (39183,-0.837518), (39184,-0.971698), (39185,-1.033887), (39186,-0.783005), (39187,-0.486132), (39188,-0.618458), (39189,-0.670422), (39190,-0.757695), (39191,-0.609461), (39192,-0.768262), (39193,-0.924276), (39194,-0.629731), (39195,-0.396495), (39196,-0.426631), (39197,-0.604479), (39198,-0.599775), (39199,-0.766008), (39200,-0.804040), (39201,-0.955872), (39202,-0.633920), (39203,-0.426237), (39204,-0.474951), (39205,-0.670909), (39206,-0.516638), (39207,-0.584400), (39208,-0.919705), (39209,-1.068756), (39210,-0.400753), (39211,-0.552584), (39212,-0.607804), (39213,-0.731302), (39214,-0.753078), (39215,-0.897477), (39216,-0.946197), (39217,-1.086413), (39218,-0.418416), (39219,-0.594869), (39220,-0.646833), (39221,-0.803310), (39222,-0.580762), (39223,-0.702400), (39224,-0.864920), (39225,-1.054378), (39226,-0.367333), (39227,-0.524274), (39228,-0.565092), (39229,-0.748977), (39230,-0.799081), (39231,-0.898891), (39232,-0.953184), (39233,-1.084577), (39234,-0.421690), (39235,-0.605105), (39236,-0.679830), (39237,-0.801474), (39238,-0.575207), (39239,-0.757695), (39240,-0.896058), (39241,-1.000050), (39242,-0.343662), (39243,-0.509432), (39244,-0.570688), (39245,-0.734129), (39246,-0.760088), (39247,-0.909133), (39248,-0.930440), (39249,-1.080881), (39250,-0.423103), (39251,-0.570752), (39252,-0.622253), (39253,-0.797315), (39254,-0.584980), (39255,-0.737744), (39256,-0.799464), (39257,-0.979629), (39258,-0.672543), (39259,-0.364529), (39260,-0.440651), (39261,-0.597128), (39262,-0.576169), (39263,-0.734500), (39264,-0.799012), (39265,-0.961989), (39266,-0.697639), (39267,-0.433282), (39268,-0.477356), (39269,-0.633833), (39270,-0.500464), (39271,-0.561257), (39272,-0.823175), (39273,-0.996841), (39274,-0.297717), (39275,-0.455122), (39276,-0.519634), (39277,-0.668216), (39278,-0.684876), (39279,-0.802801), (39280,-0.878459), (39281,-1.051192), (39282,-0.353464), (39283,-0.538745), (39284,-0.586527), (39285,-0.714207), (39286,-0.504664), (39287,-0.667648), (39288,-0.871038), (39289,-1.019156), (39290,-0.345117), (39291,-0.509954), (39292,-0.542412), (39293,-0.700286), (39294,-0.712307), (39295,-0.875284), (39296,-1.156713), (39297,-0.922087), (39298,-0.710222), (39299,-0.734778), (39300,-0.894975), (39301,-0.738382), (39302,-0.799638), (39303,-0.832097), (39304,-1.028524), (39305,-1.158057), (39306,-0.493773), (39307,-0.610308), (39308,-0.640907), (39309,-0.816426), (39310,-0.828447), (39311,-0.939872), (39312,-1.006701), (39313,-1.178507), (39314,-0.501681), (39315,-0.669774), (39316,-0.727774), (39317,-0.854064), (39318,-0.616651), (39319,-0.771733), (39320,-1.054089), (39321,-1.222182), (39322,-0.588549), (39323,-0.687895), (39324,-0.752870), (39325,-0.924213), (39326,-0.946453), (39327,-1.101534), (39328,-1.172083), (39329,-1.325774), (39330,-0.636869), (39331,-0.771049), (39332,-0.859713), (39333,-0.997612), (39334,-0.716073), (39335,-0.856758), (39336,-0.971896), (39337,-1.186432), (39338,-0.489638), (39339,-0.608489), (39340,-0.672995), (39341,-0.821113), (39342,-0.812696), (39343,-0.953845), (39344,-1.055977), (39345,-1.150214), (39346,-0.495686), (39347,-0.648907), (39348,-0.737571), (39349,-0.891262), (39350,-0.658958), (39351,-0.797321), (39352,-1.006284), (39353,-1.151616), (39354,-0.484082), (39355,-0.671217), (39356,-0.734796), (39357,-0.884304), (39358,-0.887033), (39359,-1.037474), (39360,-1.084335), (39361,-1.235703), (39362,-0.558407), (39363,-0.685161), (39364,-0.731552), (39365,-0.907077), (39366,-0.675701), (39367,-0.849830), (39368,-0.921305), (39369,-1.074063), (39370,-0.409780), (39371,-0.570903), (39372,-0.631696), (39373,-0.776095), (39374,-0.786262), (39375,-0.912546), (39376,-1.008173), (39377,-1.182302), (39378,-0.526377), (39379,-0.669386), (39380,-0.692089), (39381,-0.809550), (39382,-0.614410), (39383,-0.764382), (39384,-1.069962), (39385,-1.199502), (39386,-0.578881), (39387,-0.711201), (39388,-0.770134), (39389,-0.903387), (39390,-0.906122), (39391,-1.066312), (39392,-1.120136), (39393,-1.285443), (39394,-0.605367), (39395,-0.753948), (39396,-0.812882), (39397,-0.980042), (39398,-0.757957), (39399,-0.869376), (39400,-0.912517), (39401,-1.076427), (39402,-0.428405), (39403,-0.585809), (39404,-0.628024), (39405,-0.790538), (39406,-0.824856), (39407,-0.938134), (39408,-1.025402), (39409,-1.147046), (39410,-0.494834), (39411,-0.621118), (39412,-0.655437), (39413,-0.812377), (39414,-0.583794), (39415,-0.724009), (39416,-0.850763), (39417,-1.041611), (39418,-0.362931), (39419,-0.486892), (39420,-0.536539), (39421,-0.658640), (39422,-0.657655), (39423,-0.844327), (39424,-0.947386), (39425,-1.085748), (39426,-0.432610), (39427,-0.589094), (39428,-0.619693), (39429,-0.769202), (39430,-0.553617), (39431,-0.679444), (39432,-0.890266), (39433,-1.027232), (39434,-0.358302), (39435,-0.527322), (39436,-0.593688), (39437,-0.736697), (39438,-0.744535), (39439,-0.899159), (39440,-0.958092), (39441,-1.128965), (39442,-0.481406), (39443,-0.605367), (39444,-0.614601), (39445,-0.786871), (39446,-0.556890), (39447,-0.725910), (39448,-0.887960), (39449,-0.627786), (39450,-0.752217), (39451,-0.420509), (39452,-0.590925), (39453,-0.563460), (39454,-0.723193), (39455,-0.811387), (39456,-0.955323), (39457,-0.693295), (39458,-0.814006), (39459,-0.507846), (39460,-0.671756), (39461,-0.493798), (39462,-0.659098), (39463,-0.581007), (39464,-0.985992), (39465,-0.719781), (39466,-0.493514), (39467,-0.542228), (39468,-0.697316), (39469,-0.716299), (39470,-0.887179), (39471,-0.941929), (39472,-1.083078), (39473,-0.795503), (39474,-0.525573), (39475,-0.574750), (39476,-0.764208), (39477,-0.606688), (39478,-0.696742), (39479,-0.719914), (39480,-1.012489), (39481,-0.715616), (39482,-0.508860), (39483,-0.534819), (39484,-0.708015), (39485,-0.669874), (39486,-0.884873), (39487,-0.921051), (39488,-1.082169), (39489,-0.767649), (39490,-0.528846), (39491,-0.569664), (39492,-0.757263), (39493,-0.615534), (39494,-0.692582), (39495,-0.712036), (39496,-0.986496), (39497,-0.686378), (39498,-0.444783), (39499,-0.478631), (39500,-0.635572), (39501,-0.633661), (39502,-0.822655), (39503,-0.901563), (39504,-1.028310), (39505,-0.754204), (39506,-0.536759), (39507,-0.584084), (39508,-0.726159), (39509,-0.572822), (39510,-0.652193), (39511,-0.700444), (39512,-0.814655), (39513,-0.586992), (39514,-0.768090), (39515,-0.408981), (39516,-0.564526), (39517,-0.534280), (39518,-0.677752), (39519,-0.704632), (39520,-0.836032), (39521,-0.587003), (39522,-0.762529), (39523,-0.450796), (39524,-0.618883), (39525,-0.486910), (39526,-0.644784), (39527,-0.607100), (39528,-0.825818), (39529,-0.946066), (39530,-0.323121), (39531,-0.467063), (39532,-0.518100), (39533,-0.646244), (39534,-0.652222), (39535,-0.812419), (39536,-0.867169), (39537,-1.028757), (39538,-0.359363), (39539,-0.494476), (39540,-0.559915), (39541,-0.721965), (39542,-0.493375), (39543,-0.644743), (39544,-0.954970), (39545,-0.669718), (39546,-0.450413), (39547,-0.498201), (39548,-0.663507), (39549,-0.633719), (39550,-0.803672), (39551,-0.866781), (39552,-1.113840), (39553,-1.238728), (39554,-0.551219), (39555,-0.703057), (39556,-0.766167), (39557,-0.890597), (39558,-0.658757), (39559,-0.799443), (39560,-1.103627), (39561,-0.860177), (39562,-0.567486), (39563,-0.719324), (39564,-0.765252), (39565,-0.948667), (39566,-0.981589), (39567,-1.156182), (39568,-1.161240), (39569,-0.944258), (39570,-0.664579), (39571,-0.838245), (39572,-0.926439), (39573,-0.946819), (39574,-0.791159), (39575,-0.996872), (39576,-0.985204), (39577,-1.006981), (39578,-0.739837), (39579,-0.474090), (39580,-0.650073), (39581,-0.677422), (39582,-0.876172), (39583,-0.835702), (39584,-1.004721), (39585,-1.037643), (39586,-0.821595), (39587,-0.529374), (39588,-0.678419), (39589,-0.727133), (39590,-0.776317), (39591,-0.632729), (39592,-1.063724), (39593,-0.752455), (39594,-0.881525), (39595,-0.599986), (39596,-0.763433), (39597,-0.844201), (39598,-0.977917), (39599,-0.965317), (39600,-1.150128), (39601,-0.816104), (39602,-0.928449), (39603,-0.672458), (39604,-0.839154), (39605,-0.784751), (39606,-0.932406), (39607,-0.792074), (39608,-0.991281), (39609,-1.033496), (39610,-0.798406), (39611,-0.538695), (39612,-0.678448), (39613,-0.691865), (39614,-0.895255), (39615,-0.891020), (39616,-1.021024), (39617,-1.088780), (39618,-0.844861), (39619,-0.589333), (39620,-0.736988), (39621,-0.798244), (39622,-0.864610), (39623,-0.693157), (39624,-1.043790), (39625,-0.745063), (39626,-0.863920), (39627,-0.612106), (39628,-0.738853), (39629,-0.801042), (39630,-0.972385), (39631,-0.962571), (39632,-1.096287), (39633,-0.783628), (39634,-0.947538), (39635,-0.701296), (39636,-0.855920), (39637,-0.813590), (39638,-0.961708), (39639,-0.788396), (39640,-0.948593), (39641,-0.987551), (39642,-0.771040), (39643,-0.489037), (39644,-0.624607), (39645,-0.685870), (39646,-0.866035), (39647,-0.871550), (39648,-1.016882), (39649,-1.045621), (39650,-0.798922), (39651,-0.576368), (39652,-0.719840), (39653,-0.762518), (39654,-0.831207), (39655,-0.670900), (39656,-0.845956), (39657,-0.869592), (39658,-0.658190), (39659,-0.396620), (39660,-0.563316), (39661,-0.588806), (39662,-0.766185), (39663,-0.776815), (39664,-0.942579), (39665,-1.024273), (39666,-0.752490), (39667,-0.474664), (39668,-0.604668), (39669,-0.666387), (39670,-0.736472), (39671,-0.583592), (39672,-0.759581), (39673,-0.796686), (39674,-0.555553), (39675,-0.303739), (39676,-0.470435), (39677,-0.529375), (39678,-0.678883), (39679,-0.662106), (39680,-0.836699), (39681,-0.908638), (39682,-0.665188), (39683,-0.385966), (39684,-0.563815), (39685,-0.589768), (39686,-0.645451), (39687,-0.499540), (39688,-0.828345), (39689,-0.881705), (39690,-0.666590), (39691,-0.395734), (39692,-0.538273), (39693,-0.587920), (39694,-0.779701), (39695,-0.734584), (39696,-0.907786), (39697,-0.938385), (39698,-0.687967), (39699,-0.426866), (39700,-0.618640), (39701,-0.646453), (39702,-0.710966), (39703,-0.563664), (39704,-0.908261), (39705,-1.065666), (39706,-0.402315), (39707,-0.594089), (39708,-0.650706), (39709,-0.763521), (39710,-0.765786), (39711,-0.932946), (39712,-1.004884), (39713,-1.176227), (39714,-0.514730), (39715,-0.670744), (39716,-0.732000), (39717,-0.877332), (39718,-0.645022), (39719,-0.757844), (39720,-0.873445), (39721,-1.040141), (39722,-0.365639), (39723,-0.511897), (39724,-0.559685), (39725,-0.698510), (39726,-0.692416), (39727,-0.823809), (39728,-0.889249), (39729,-1.021105), (39730,-0.333134), (39731,-0.514695), (39732,-0.587561), (39733,-0.733356), (39734,-0.455993), (39735,-0.597612), (39736,-0.775454), (39737,-0.933328), (39738,-0.282050), (39739,-0.445027), (39740,-0.495601), (39741,-0.645116), (39742,-0.669672), (39743,-0.834515), (39744,-0.890192), (39745,-1.043420), (39746,-0.390289), (39747,-0.525858), (39748,-0.596870), (39749,-0.774719), (39750,-0.545665), (39751,-0.682631), (39752,-0.852114), (39753,-0.985367), (39754,-0.291823), (39755,-0.464556), (39756,-0.556933), (39757,-0.666961), (39758,-0.715212), (39759,-0.835459), (39760,-0.861419), (39761,-1.000244), (39762,-0.349893), (39763,-0.501731), (39764,-0.569486), (39765,-0.716208), (39766,-0.481582), (39767,-0.643169), (39768,-0.891618), (39769,-1.017438), (39770,-0.379165), (39771,-0.531467), (39772,-0.585754), (39773,-0.727366), (39774,-0.744033), (39775,-0.846165), (39776,-0.930183), (39777,-1.089447), (39778,-0.418194), (39779,-0.557953), (39780,-0.608527), (39781,-0.744566), (39782,-0.529914), (39783,-0.658984), (39784,-0.949700), (39785,-0.658405), (39786,-0.351318), (39787,-0.517552), (39788,-0.571839), (39789,-0.754327), (39790,-0.740800), (39791,-0.895424), (39792,-0.981295), (39793,-0.709975), (39794,-0.452124), (39795,-0.636936), (39796,-0.680077), (39797,-0.764558), (39798,-0.594032), (39799,-0.804855), (39800,-0.865648), (39801,-1.027235), (39802,-0.351805), (39803,-0.471589), (39804,-0.554674), (39805,-0.698609), (39806,-0.694838), (39807,-0.833201), (39808,-1.178731), (39809,-1.224658), (39810,-0.990958), (39811,-0.703377), (39812,-0.863111), (39813,-0.923434), (39814,-0.998165), (39815,-0.856900), (39816,-1.069119), (39817,-1.151740), (39818,-0.914791), (39819,-0.642538), (39820,-0.753499), (39821,-0.813822), (39822,-0.973556), (39823,-0.963742), (39824,-1.063088), (39825,-1.148966), (39826,-0.922235), (39827,-0.616075), (39828,-0.764657), (39829,-0.831023), (39830,-0.933618), (39831,-0.770989), (39832,-1.020828), (39833,-1.092773), (39834,-0.870682), (39835,-0.582174), (39836,-0.722859), (39837,-0.787835), (39838,-0.968927), (39839,-0.960046), (39840,-1.110024), (39841,-1.167561), (39842,-0.924575), (39843,-0.629568), (39844,-0.818556), (39845,-0.849155), (39846,-0.928532), (39847,-0.826747), (39848,-0.862919), (39849,-1.031939), (39850,-0.671904), (39851,-0.814443), (39852,-0.555665), (39853,-0.742800), (39854,-0.801269), (39855,-0.926163), (39856,-0.920995), (39857,-1.083046), (39858,-0.755058), (39859,-0.868336), (39860,-0.606766), (39861,-0.784151), (39862,-0.745540), (39863,-0.901091), (39864,-1.018082), (39865,-1.175956), (39866,-0.832639), (39867,-0.993757), (39868,-0.733589), (39869,-0.860336), (39870,-0.943890), (39871,-1.080393), (39872,-1.084518), (39873,-1.209875), (39874,-0.876307), (39875,-1.022102), (39876,-0.787939), (39877,-0.940704), (39878,-0.899769), (39879,-1.019554), (39880,-0.924738), (39881,-1.109556), (39882,-0.754623), (39883,-0.882304), (39884,-0.611447), (39885,-0.754913), (39886,-0.853332), (39887,-1.009346), (39888,-0.999069), (39889,-1.127213), (39890,-0.784359), (39891,-0.938514), (39892,-0.693668), (39893,-0.819489), (39894,-0.782274), (39895,-0.938288), (39896,-0.981893), (39897,-1.121652), (39898,-0.817815), (39899,-0.960823), (39900,-0.680211), (39901,-0.867809), (39902,-0.894226), (39903,-1.041417), (39904,-1.051115), (39905,-1.212238), (39906,-0.864276), (39907,-1.022143), (39908,-0.731312), (39909,-0.910551), (39910,-0.856611), (39911,-0.999620), (39912,-0.855105), (39913,-0.995790), (39914,-0.678485), (39915,-0.849827), (39916,-0.564106), (39917,-0.720583), (39918,-0.775340), (39919,-0.949932), (39920,-0.922930), (39921,-1.088700), (39922,-0.722622), (39923,-0.871204), (39924,-0.612890), (39925,-0.779586), (39926,-0.766523), (39927,-0.904422), (39928,-0.651217), (39929,-0.778891), (39930,-0.852689), (39931,-0.608777), (39932,-0.332341), (39933,-0.461881), (39934,-0.544502), (39935,-0.741392), (39936,-0.717183), (39937,-0.870411), (39938,-0.931204), (39939,-0.671029), (39940,-0.402959), (39941,-0.531566), (39942,-0.589573), (39943,-0.666157), (39944,-0.680965), (39945,-0.854161), (39946,-0.907984), (39947,-0.711448), (39948,-0.410397), (39949,-0.532968), (39950,-0.637887), (39951,-0.783682), (39952,-0.797562), (39953,-0.926633), (39954,-0.983706), (39955,-0.752336), (39956,-0.467077), (39957,-0.621695), (39958,-0.660660), (39959,-0.706124), (39960,-0.766911), (39961,-0.830027), (39962,-1.005083), (39963,-0.311538), (39964,-0.426213), (39965,-0.516267), (39966,-0.692255), (39967,-0.730751), (39968,-0.866327), (39969,-0.971709), (39970,-1.104499), (39971,-0.428599), (39972,-0.593443), (39973,-0.630541), (39974,-0.773550), (39975,-0.539387), (39976,-0.981998), (39977,-1.059046), (39978,-0.781683), (39979,-0.516400), (39980,-0.688669), (39981,-0.742963), (39982,-0.906873), (39983,-0.880340), (39984,-1.034958), (39985,-1.113866), (39986,-0.849972), (39987,-0.574939), (39988,-0.733740), (39989,-0.735072), (39990,-0.815376), (39991,-0.670398), (39992,-0.751160), (39993,-0.823098), (39994,-1.035317), (39995,-0.344096), (39996,-0.486635), (39997,-0.512124), (39998,-0.662566), (39999,-0.685732), (40000,-0.836174), (40001,-0.885821), (40002,-1.021860), (40003,-0.380338), (40004,-0.558643), (40005,-0.594352), (40006,-0.717849), (40007,-0.496228), (40008,-0.697765), (40009,-0.758094), (40010,-0.889488), (40011,-0.240996), (40012,-0.409089), (40013,-0.487997), (40014,-0.619853), (40015,-0.611436), (40016,-0.779529), (40017,-0.886765), (40018,-1.020018), (40019,-0.365026), (40020,-0.529863), (40021,-0.571151), (40022,-0.711367), (40023,-0.499038), (40024,-0.757243), (40025,-0.797598), (40026,-0.954075), (40027,-0.267494), (40028,-0.415142), (40029,-0.451784), (40030,-0.620804), (40031,-0.641184), (40032,-0.766077), (40033,-0.803176), (40034,-0.987524), (40035,-0.306985), (40036,-0.454171), (40037,-0.523792), (40038,-0.717890), (40039,-0.462825), (40040,-0.823221), (40041,-0.853356), (40042,-0.630339), (40043,-0.286096), (40044,-0.469511), (40045,-0.540523), (40046,-0.693751), (40047,-0.689510), (40048,-0.848310), (40049,-0.920249), (40050,-0.670764), (40051,-0.404547), (40052,-0.558701), (40053,-0.636683), (40054,-0.686793), (40055,-0.529273), (40056,-0.951439), (40057,-0.995507), (40058,-0.731157), (40059,-0.504426), (40060,-0.653008), (40061,-0.705441), (40062,-0.880497), (40063,-0.857215), (40064,-1.233865), (40065,-1.294652), (40066,-1.062348), (40067,-0.748762), (40068,-0.890838), (40069,-0.972532), (40070,-1.043081), (40071,-0.870232), (40072,-1.102419), (40073,-1.140451), (40074,-0.929982), (40075,-0.627999), (40076,-0.802128), (40077,-0.839696), (40078,-1.059811), (40079,-1.046748), (40080,-1.187433), (40081,-1.239397), (40082,-0.960645), (40083,-0.719055), (40084,-0.837906), (40085,-0.870365), (40086,-0.953450), (40087,-0.831696), (40088,-0.964949), (40089,-0.979293), (40090,-1.133911), (40091,-0.503070), (40092,-0.663731), (40093,-0.712445), (40094,-0.884714), (40095,-0.880480), (40096,-1.035098), (40097,-1.054551), (40098,-1.237503), (40099,-0.554178), (40100,-0.691144), (40101,-0.751010), (40102,-0.922816), (40103,-0.693762), (40104,-0.917590), (40105,-1.062459), (40106,-0.752116), (40107,-0.872364), (40108,-0.611726), (40109,-0.744052), (40110,-0.821564), (40111,-0.984547), (40112,-0.974734), (40113,-1.120065), (40114,-0.774426), (40115,-0.919758), (40116,-0.647968), (40117,-0.802586), (40118,-0.763511), (40119,-0.929281), (40120,-1.051388), (40121,-1.190678), (40122,-0.823673), (40123,-0.985260), (40124,-0.716727), (40125,-0.854619), (40126,-0.941423), (40127,-1.096974), (40128,-1.079734), (40129,-1.270582), (40130,-0.921223), (40131,-1.084206), (40132,-0.822172), (40133,-0.970754), (40134,-0.922393), (40135,-1.071902), (40136,-0.965013), (40137,-1.096407), (40138,-0.799076), (40139,-0.926286), (40140,-0.648467), (40141,-0.817017), (40142,-0.893138), (40143,-1.055189), (40144,-1.029589), (40145,-1.193963), (40146,-0.875724), (40147,-1.013623), (40148,-0.756699), (40149,-0.864404), (40150,-0.841591), (40151,-1.020830), (40152,-0.872596), (40153,-1.045335), (40154,-1.106591), (40155,-0.821796), (40156,-0.554189), (40157,-0.720422), (40158,-0.740339), (40159,-0.943266), (40160,-0.980371), (40161,-1.109441), (40162,-1.135864), (40163,-0.922602), (40164,-0.623411), (40165,-0.796144), (40166,-0.846718), (40167,-0.921913), (40168,-0.787154), (40169,-0.932479), (40170,-0.981663), (40171,-0.722879), (40172,-0.450163), (40173,-0.617792), (40174,-0.657214), (40175,-0.826697), (40176,-0.797378), (40177,-0.953856), (40178,-0.990961), (40179,-0.774449), (40180,-0.488727), (40181,-0.622907), (40182,-0.643294), (40183,-0.731024), (40184,-0.619490), (40185,-0.808484), (40186,-0.866948), (40187,-0.629071), (40188,-0.368897), (40189,-0.518412), (40190,-0.564339), (40191,-0.739395), (40192,-0.743983), (40193,-0.906497), (40194,-0.956608), (40195,-0.728487), (40196,-0.443229), (40197,-0.620144), (40198,-0.672108), (40199,-0.740797), (40200,-0.737489), (40201,-0.879102), (40202,-0.925962), (40203,-0.669501), (40204,-0.391212), (40205,-0.547690), (40206,-0.575502), (40207,-0.801190), (40208,-0.805778), (40209,-0.959006), (40210,-0.982642), (40211,-0.723395), (40212,-0.467867), (40213,-0.593224), (40214,-0.655870), (40215,-0.728742), (40216,-0.812759), (40217,-0.898637), (40218,-1.027243), (40219,-0.342985), (40220,-0.486457), (40221,-0.547713), (40222,-0.688862), (40223,-0.699487), (40224,-0.903810), (40225,-0.997119), (40226,-1.085313), (40227,-0.435431), (40228,-0.596085), (40229,-0.629941), (40230,-0.835654), (40231,-0.604740), (40232,-0.853189), (40233,-0.910269), (40234,-1.078819), (40235,-0.421505), (40236,-0.562654), (40237,-0.592789), (40238,-0.753450), (40239,-0.773830), (40240,-0.890821), (40241,-0.945115), (40242,-1.096946), (40243,-0.454027), (40244,-0.614224), (40245,-0.653646), (40246,-0.812910), (40247,-0.573174), (40248,-0.804441), (40249,-0.879629), (40250,-1.004523), (40251,-0.346739), (40252,-0.510186), (40253,-0.594203), (40254,-0.733029), (40255,-0.754342), (40256,-0.879229), (40257,-0.927017), (40258,-1.098360), (40259,-0.384840), (40260,-0.552927), (40261,-0.559838), (40262,-0.732577), (40263,-0.490518), (40264,-0.735711), (40265,-0.798364), (40266,-0.959024), (40267,-0.294740), (40268,-0.421024), (40269,-0.439544), (40270,-0.617856), (40271,-0.655888), (40272,-0.824445), (40273,-0.861080), (40274,-0.975755), (40275,-0.304965), (40276,-0.501855), (40277,-0.544070), (40278,-0.720522), (40279,-0.511437), (40280,-0.790543), (40281,-0.842044), (40282,-0.962761), (40283,-0.314732), (40284,-0.484679), (40285,-0.517601), (40286,-0.671755), (40287,-0.690745), (40288,-0.876020), (40289,-0.926131), (40290,-1.107693), (40291,-0.413215), (40292,-0.554827), (40293,-0.609114), (40294,-0.747947), (40295,-0.547690), (40296,-0.913659), (40297,-0.977232), (40298,-0.716594), (40299,-0.426696), (40300,-0.597106), (40301,-0.655112), (40302,-0.809730), (40303,-0.833366), (40304,-0.961046), (40305,-1.029735), (40306,-0.794175), (40307,-0.467577), (40308,-0.643566), (40309,-0.703896), (40310,-0.732172), (40311,-0.618314), (40312,-1.045590), (40313,-1.104524), (40314,-0.864788), (40315,-0.530300), (40316,-0.665406), (40317,-0.728059), (40318,-0.936095), (40319,-0.929538), (40320,-1.051175), (40321,-1.109645), (40322,-1.286561), (40323,-0.612058), (40324,-0.738341), (40325,-0.805177), (40326,-0.953289), (40327,-0.724705), (40328,-0.977794), (40329,-1.058561), (40330,-1.218758), (40331,-0.521494), (40332,-0.709556), (40333,-0.756880), (40334,-0.884554), (40335,-0.864064), (40336,-1.012182), (40337,-1.094340), (40338,-1.248031), (40339,-0.554943), (40340,-0.711421), (40341,-0.801011), (40342,-0.949593), (40343,-0.694535), (40344,-0.930435), (40345,-0.982869), (40346,-1.149102), (40347,-0.497360), (40348,-0.606456), (40349,-0.712308), (40350,-0.852060), (40351,-0.859435), (40352,-0.967610), (40353,-1.036299), (40354,-1.191380), (40355,-0.523383), (40356,-0.638051), (40357,-0.716496), (40358,-0.877620), (40359,-0.671327), (40360,-1.008492), (40361,-1.176121), (40362,-0.836054), (40363,-0.980453), (40364,-0.688695), (40365,-0.860501), (40366,-0.949628), (40367,-1.110282), (40368,-1.076317), (40369,-1.227685), (40370,-0.897838), (40371,-1.028304), (40372,-0.762557), (40373,-0.930650), (40374,-0.863705), (40375,-1.005317), (40376,-0.898892), (40377,-1.039578), (40378,-1.110590), (40379,-0.839733), (40380,-0.563304), (40381,-0.734177), (40382,-0.764313), (40383,-0.974672), (40384,-0.989016), (40385,-1.134811), (40386,-1.184921), (40387,-0.918241), (40388,-0.664103), (40389,-0.808508), (40390,-0.854436), (40391,-0.935204), (40392,-0.777214), (40393,-0.968068), (40394,-1.032574), (40395,-0.794698), (40396,-0.512689), (40397,-0.690074), (40398,-0.714631), (40399,-0.875755), (40400,-0.891025), (40401,-1.053545), (40402,-1.127807), (40403,-0.853694), (40404,-0.563333), (40405,-0.714701), (40406,-0.756909), (40407,-0.827458), (40408,-0.863630), (40409,-1.027076), (40410,-1.071151), (40411,-0.804934), (40412,-0.514572), (40413,-0.690092), (40414,-0.724410), (40415,-0.921294), (40416,-0.910554), (40417,-1.061458), (40418,-1.116678), (40419,-0.886698), (40420,-0.613518), (40421,-0.784391), (40422,-0.815460), (40423,-0.905514), (40424,-0.763786), (40425,-0.930019), (40426,-0.971764), (40427,-0.736674), (40428,-0.453275), (40429,-0.610686), (40430,-0.656613), (40431,-0.854894), (40432,-0.797241), (40433,-0.931421), (40434,-1.044236), (40435,-0.819365), (40436,-0.508559), (40437,-0.665036), (40438,-0.723976), (40439,-0.803810), (40440,-0.766126), (40441,-0.904958), (40442,-0.963891), (40443,-0.739484), (40444,-0.450512), (40445,-0.591661), (40446,-0.667783), (40447,-0.858167), (40448,-0.826525), (40449,-0.989039), (40450,-1.016388), (40451,-0.774329), (40452,-0.534130), (40453,-0.632543), (40454,-0.706341), (40455,-0.769457), (40456,-0.785191), (40457,-0.937492), (40458,-1.028009), (40459,-0.792456), (40460,-0.509057), (40461,-0.659499), (40462,-0.705890), (40463,-0.877232), (40464,-0.840481), (40465,-1.040621), (40466,-1.068434), (40467,-0.823119), (40468,-0.511386), (40469,-0.681339), (40470,-0.697999), (40471,-0.785273), (40472,-0.720187), (40473,-0.767042), (40474,-0.917946), (40475,-0.677747), (40476,-0.436615), (40477,-0.486725), (40478,-0.662708), (40479,-0.654290), (40480,-0.838639), (40481,-0.872030), (40482,-1.010856), (40483,-0.757645), (40484,-0.500264), (40485,-0.561520), (40486,-0.755618), (40487,-0.635724), (40488,-0.890209), (40489,-0.938460), (40490,-1.084255), (40491,-0.400929), (40492,-0.573199), (40493,-0.623303), (40494,-0.793256), (40495,-0.801557), (40496,-0.942706), (40497,-0.996530), (40498,-1.149294), (40499,-0.489657), (40500,-0.616404), (40501,-0.679056), (40502,-0.797907), (40503,-0.564677), (40504,-0.922280), (40505,-0.997475), (40506,-1.132118), (40507,-0.488735), (40508,-0.625708), (40509,-0.662806), (40510,-0.816034), (40511,-0.817836), (40512,-0.994288), (40513,-1.056008), (40514,-1.192511), (40515,-0.553775), (40516,-0.700496), (40517,-0.733419), (40518,-0.879214), (40519,-0.640874), (40520,-0.917657), (40521,-0.970084), (40522,-1.113093), (40523,-0.412579), (40524,-0.585782), (40525,-0.665153), (40526,-0.808625), (40527,-0.825286), (40528,-0.947856), (40529,-1.030014), (40530,-1.182315), (40531,-0.479942), (40532,-0.640132), (40533,-0.696749), (40534,-0.846257), (40535,-0.600948), (40536,-0.698434), (40537,-0.761550), (40538,-0.911522), (40539,-0.657854), (40540,-0.412081), (40541,-0.436175), (40542,-0.548990), (40543,-0.545682), (40544,-0.752328), (40545,-0.809865), (40546,-0.971915), (40547,-0.694559), (40548,-0.473865), (40549,-0.503074), (40550,-0.647936), (40551,-0.527579), (40552,-0.952068), (40553,-0.991027), (40554,-0.751291), (40555,-0.465105), (40556,-0.619266), (40557,-0.672626), (40558,-0.823061), (40559,-0.839265), (40560,-1.007352), (40561,-1.011940), (40562,-0.794965), (40563,-0.505530), (40564,-0.665257), (40565,-0.692143), (40566,-0.763619), (40567,-0.599592), (40568,-0.814135), (40569,-0.865635), (40570,-1.015150), (40571,-0.366658), (40572,-0.537531), (40573,-0.617372), (40574,-0.758984), (40575,-0.754743), (40576,-1.053361), (40577,-1.194973), (40578,-0.881844), (40579,-1.034609), (40580,-0.768861), (40581,-0.892822), (40582,-0.858394), (40583,-1.028340), (40584,-0.992058), (40585,-1.107660), (40586,-0.788031), (40587,-0.919888), (40588,-0.618374), (40589,-0.780894), (40590,-0.876521), (40591,-1.044144), (40592,-1.077536), (40593,-1.207996), (40594,-0.868399), (40595,-1.017444), (40596,-0.738222), (40597,-0.907241), (40598,-0.922048), (40599,-1.032077), (40600,-0.888958), (40601,-1.021285), (40602,-1.057920), (40603,-0.830263), (40604,-0.566369), (40605,-0.715420), (40606,-0.785036), (40607,-0.972634), (40608,-0.963753), (40609,-1.131377), (40610,-1.210748), (40611,-0.930136), (40612,-0.608184), (40613,-0.802751), (40614,-0.845892), (40615,-0.893216), (40616,-0.919633), (40617,-1.044526), (40618,-0.716538), (40619,-0.912032), (40620,-0.588221), (40621,-0.739126), (40622,-0.838008), (40623,-0.995882), (40624,-0.957734), (40625,-1.108639), (40626,-0.734665), (40627,-0.897179), (40628,-0.653730), (40629,-0.794415), (40630,-0.733970), (40631,-0.905776), (40632,-1.050644), (40633,-1.201079), (40634,-0.863805), (40635,-0.985443), (40636,-0.706227), (40637,-0.876173), (40638,-0.962977), (40639,-1.118991), (40640,-1.111501), (40641,-1.269375), (40642,-0.922338), (40643,-1.097394), (40644,-0.835367), (40645,-0.994167), (40646,-0.969952), (40647,-1.112034), (40648,-0.953117), (40649,-1.111918), (40650,-0.754669), (40651,-0.924152), (40652,-0.656082), (40653,-0.782829), (40654,-0.855701), (40655,-1.003349), (40656,-1.022339), (40657,-1.156056), (40658,-0.816922), (40659,-0.973863), (40660,-0.684891), (40661,-0.808388), (40662,-0.808794), (40663,-0.908140), (40664,-0.844451), (40665,-1.020897), (40666,-1.060788), (40667,-0.807583), (40668,-0.546013), (40669,-0.680199), (40670,-0.727516), (40671,-0.909542), (40672,-0.952683), (40673,-1.103587), (40674,-1.163454), (40675,-0.917675), (40676,-0.628240), (40677,-0.813052), (40678,-0.817177), (40679,-0.890975), (40680,-0.694902), (40681,-0.764054), (40682,-0.921458), (40683,-0.634346), (40684,-0.770386), (40685,-0.466549), (40686,-0.633245), (40687,-0.724695), (40688,-0.879313), (40689,-0.863933), (40690,-1.010655), (40691,-0.697989), (40692,-0.861436), (40693,-0.573861), (40694,-0.711753), (40695,-0.681045), (40696,-0.661475), (40697,-0.825849), (40698,-0.923805), (40699,-0.675240), (40700,-0.406243), (40701,-0.563647), (40702,-0.593783), (40703,-0.768375), (40704,-0.700040), (40705,-0.896467), (40706,-0.919634), (40707,-0.698939), (40708,-0.408108), (40709,-0.596639), (40710,-0.662078), (40711,-0.709859), (40712,-0.677754), (40713,-0.754339), (40714,-0.905244), (40715,-0.575396), (40716,-0.694717), (40717,-0.428969), (40718,-0.591483), (40719,-0.646703), (40720,-0.807357), (40721,-0.803123), (40722,-0.963313), (40723,-0.613497), (40724,-0.777871), (40725,-0.524660), (40726,-0.681607), (40727,-0.648568), (40728,-0.793900), (40729,-0.830999), (40730,-0.977264), (40731,-0.265135), (40732,-0.466201), (40733,-0.519098), (40734,-0.690905), (40735,-0.724753), (40736,-0.866835), (40737,-0.890929), (40738,-1.058095), (40739,-0.413780), (40740,-0.527064), (40741,-0.619904), (40742,-0.800070), (40743,-0.551048), (40744,-0.699160), (40745,-0.876545), (40746,-0.903425), (40747,-0.689699), (40748,-0.391905), (40749,-0.577180), (40750,-0.612889), (40751,-0.767513), (40752,-0.741907), (40753,-0.922536), (40754,-1.007480), (40755,-0.737093), (40756,-0.476919), (40757,-0.612959), (40758,-0.693257), (40759,-0.777737), (40760,-0.822738), (40761,-0.855661), (40762,-1.018644), (40763,-0.354360), (40764,-0.496899), (40765,-0.564662), (40766,-0.714170), (40767,-0.722477), (40768,-0.877559), (40769,-0.937888), (40770,-1.062312), (40771,-0.410107), (40772,-0.562872), (40773,-0.635274), (40774,-0.755521), (40775,-0.493951), (40776,-0.660184), (40777,-0.858001), (40778,-0.876991), (40779,-0.648870), (40780,-0.333418), (40781,-0.457379), (40782,-0.539073), (40783,-0.756402), (40784,-0.716864), (40785,-0.901675), (40786,-0.920202), (40787,-0.703221), (40788,-0.402177), (40789,-0.585129), (40790,-0.635239), (40791,-0.707178), (40792,-0.721052), (40793,-0.775345), (40794,-0.936469), (40795,-0.273575), (40796,-0.410078), (40797,-0.482487), (40798,-0.626422), (40799,-0.645875), (40800,-0.781915), (40801,-0.863146), (40802,-1.026586), (40803,-0.353943), (40804,-0.506708), (40805,-0.565177), (40806,-0.709576), (40807,-0.504210), (40808,-0.778670), (40809,-0.933758), (40810,-0.589508), (40811,-0.713006), (40812,-0.447258), (40813,-0.595840), (40814,-0.694723), (40815,-0.850274), (40816,-0.810266), (40817,-0.982536), (40818,-0.642938), (40819,-0.801739), (40820,-0.494646), (40821,-0.650660), (40822,-0.627847), (40823,-0.761564), (40824,-0.881348), (40825,-1.061513), (40826,-0.740488), (40827,-0.868632), (40828,-0.578270), (40829,-0.706877), (40830,-0.812259), (40831,-0.967810), (40832,-0.763377), (40833,-0.512026), (40834,-0.563990), (40835,-0.717217), (40836,-0.416167), (40837,-0.509477), (40838,-0.578166), (40839,-0.723497), (40840,-0.648187), (40841,-0.403811), (40842,-0.462281), (40843,-0.620148), (40844,-0.381808), (40845,-0.547572), (40846,-0.616261), (40847,-0.762989), (40848,-0.728091), (40849,-0.479532), (40850,-0.524064), (40851,-0.702376), (40852,-0.415727), (40853,-0.501598), (40854,-0.524771), (40855,-0.683572), (40856,-0.499107), (40857,-0.636073), (40858,-0.322024), (40859,-0.473855), (40860,-0.205322), (40861,-0.390133), (40862,-0.451853), (40863,-0.581856), (40864,-0.590621), (40865,-0.752208), (40866,-0.374058), (40867,-0.555150), (40868,-0.286153), (40869,-0.435198), (40870,-0.397520), (40871,-0.529840), (40872,-0.649160), (40873,-0.298875), (40874,-0.455352), (40875,-0.546339), (40876,-0.673086), (40877,-0.448678), (40878,-0.594010), (40879,-0.644114), (40880,-0.797805), (40881,-0.398284), (40882,-0.523178), (40883,-0.580721), (40884,-0.702358), (40885,-0.337207), (40886,-0.515056), (40887,-0.569343), (40888,-0.673799), (40889,-0.365779), (40890,-0.508788), (40891,-0.547283), (40892,-0.714449), (40893,-0.473317), (40894,-0.652555), (40895,-0.672935), (40896,-0.825230), (40897,-0.403880), (40898,-0.578010), (40899,-0.628120), (40900,-0.800390), (40901,-0.437562), (40902,-0.565705), (40903,-0.618139), (40904,-0.583241), (40905,-0.262222), (40906,-0.434955), (40907,-0.505967), (40908,-0.655938), (40909,-0.387405), (40910,-0.570826), (40911,-0.645088), (40912,-0.776018), (40913,-0.353735), (40914,-0.483739), (40915,-0.545458), (40916,-0.707509), (40917,-0.348400), (40918,-0.491403), (40919,-0.602827), (40920,-0.543315), (40921,-0.605967), (40922,-0.347183), (40923,-0.401007), (40924,-0.565850), (40925,-0.268983), (40926,-0.423600), (40927,-0.481607), (40928,-0.650157), (40929,-0.627344), (40930,-0.380639), (40931,-0.467906), (40932,-0.605342), (40933,-0.343308), (40934,-0.428252), (40935,-0.463967), (40936,-0.420710), (40937,-0.475460), (40938,-0.245480), (40939,-0.289084), (40940,-0.425130), (40941,-0.150554), (40942,-0.353944), (40943,-0.402195), (40944,-0.567965), (40945,-0.535390), (40946,-0.298446), (40947,-0.356916), (40948,-0.486913), (40949,-0.221629), (40950,-0.347920), (40951,-0.421718), (40952,-0.368242), (40953,-0.428101), (40954,-0.160501), (40955,-0.236153), (40956,-0.396350), (40957,-0.125493), (40958,-0.280111), (40959,-0.325575), (40960,-0.489486), (40961,-0.498720), (40962,-0.254338), (40963,-0.323027), (40964,-0.458139), (40965,-0.194246), (40966,-0.247606), (40967,-0.326514), (40968,-0.391953), (40969,-0.471788), (40970,-0.237624), (40971,-0.324428), (40972,-0.448389), (40973,-0.200294), (40974,-0.355844), (40975,-0.406418), (40976,-0.545244), (40977,-0.540077), (40978,-0.260397), (40979,-0.325830), (40980,-0.487887), (40981,-0.220744), (40982,-0.302901), (40983,-0.373913), (40984,-0.529927), (40985,-0.685009), (40986,-0.336582), (40987,-0.463336), (40988,-0.184114), (40989,-0.328982), (40990,-0.394885), (40991,-0.571800), (40992,-0.542945), (40993,-0.687343), (40994,-0.383970), (40995,-0.505614), (40996,-0.238007), (40997,-0.409350), (40998,-0.380494), (40999,-0.513747), (41000,-0.413359), (41001,-0.596310), (41002,-0.226520), (41003,-0.365345), (41004,-0.082873), (41005,-0.224492), (41006,-0.308509), (41007,-0.492851), (41008,-0.492800), (41009,-0.625120), (41010,-0.299455), (41011,-0.464755), (41012,-0.126084), (41013,-0.261661), (41014,-0.252310), (41015,-0.438981), (41016,-0.410589), (41017,-0.568463), (41018,-0.210745), (41019,-0.378368), (41020,-0.129346), (41021,-0.283037), (41022,-0.337324), (41023,-0.479869), (41024,-0.476562), (41025,-0.626070), (41026,-0.274857), (41027,-0.416470), (41028,-0.137254), (41029,-0.303487), (41030,-0.256517), (41031,-0.416244), (41032,-0.364627), (41033,-0.518318), (41034,-0.185221), (41035,-0.344021), (41036,-0.108925), (41037,-0.262153), (41038,-0.304831), (41039,-0.430188), (41040,-0.445922), (41041,-0.581961), (41042,-0.230285), (41043,-0.420670), (41044,-0.148423), (41045,-0.326265), (41046,-0.259784), (41047,-0.426943), (41048,-0.488669), (41049,-0.637714), (41050,-0.278599), (41051,-0.481996), (41052,-0.149825), (41053,-0.300730), (41054,-0.364772), (41055,-0.534719), (41056,-0.525838), (41057,-0.675810), (41058,-0.311591), (41059,-0.455064), (41060,-0.167482), (41061,-0.318387), (41062,-0.302073), (41063,-0.447868), (41064,-0.497516), (41065,-0.245237), (41066,-0.290232), (41067,-0.416522), (41068,-0.160061), (41069,-0.352769), (41070,-0.405202), (41071,-0.573295), (41072,-0.555122), (41073,-0.315850), (41074,-0.350162), (41075,-0.530334), (41076,-0.258081), (41077,-0.344421), (41078,-0.380130), (41079,-0.552863), (41080,-0.552341), (41081,-0.283344), (41082,-0.363179), (41083,-0.515480), (41084,-0.237654), (41085,-0.433612), (41086,-0.510196), (41087,-0.654602), (41088,-0.614594), (41089,-0.709294), (41090,-0.464918), (41091,-0.320867), (41092,-0.458766), (41093,-0.495401), (41094,-0.562694), (41095,-0.270472), (41096,-0.431596), (41097,-0.579714), (41098,-0.245684), (41099,-0.444897), (41100,-0.436010), (41101,-0.572982), (41102,-0.600332), (41103,-0.785143), (41104,-0.485953), (41105,-0.638711), (41106,-0.317692), (41107,-0.479742), (41108,-0.353343), (41109,-0.472663), (41110,-0.477715), (41111,-0.636979), (41112,-0.473422), (41113,-0.625254), (41114,-0.296333), (41115,-0.437018), (41116,-0.434637), (41117,-0.586938), (41118,-0.657487), (41119,-0.772155), (41120,-0.509658), (41121,-0.667068), (41122,-0.338611), (41123,-0.460718), (41124,-0.339428), (41125,-0.526562), (41126,-0.519541), (41127,-0.662080), (41128,-0.626262), (41129,-0.371197), (41130,-0.444526), (41131,-0.577779), (41132,-0.594909), (41133,-0.784831), (41134,-0.834478), (41135,-0.987705), (41136,-0.690368), (41137,-0.476180), (41138,-0.527217), (41139,-0.682768), (41140,-0.535003), (41141,-0.594400), (41142,-0.618963), (41143,-0.775904), (41144,-0.509230), (41145,-0.698681), (41146,-0.358614), (41147,-0.482581), (41148,-0.484383), (41149,-0.587442), (41150,-0.705367), (41151,-0.869740), (41152,-0.593311), (41153,-0.736319), (41154,-0.385570), (41155,-0.512317), (41156,-0.384058), (41157,-0.530786), (41158,-0.502857), (41159,-0.641683), (41160,-0.394984), (41161,-0.566321), (41162,-0.237869), (41163,-0.383201), (41164,-0.391966), (41165,-0.542870), (41166,-0.653832), (41167,-0.808913), (41168,-0.521801), (41169,-0.652731), (41170,-0.324736), (41171,-0.436625), (41172,-0.306975), (41173,-0.410034), (41174,-0.396044), (41175,-0.532547), (41176,-0.421945), (41177,-0.599788), (41178,-0.245782), (41179,-0.404120), (41180,-0.402208), (41181,-0.554039), (41182,-0.650136), (41183,-0.781992), (41184,-0.448431), (41185,-0.603513), (41186,-0.284811), (41187,-0.459403), (41188,-0.331613), (41189,-0.445355), (41190,-0.433224), (41191,-0.563691), (41192,-0.285402), (41193,-0.436770), (41194,-0.095776), (41195,-0.220664), (41196,-0.246623), (41197,-0.359901), (41198,-0.453674), (41199,-0.634766), (41200,-0.356477), (41201,-0.513424), (41202,-0.152919), (41203,-0.302891), (41204,-0.192753), (41205,-0.376631), (41206,-0.306900), (41207,-0.467097), (41208,-0.335587), (41209,-0.480450), (41210,-0.109732), (41211,-0.268996), (41212,-0.248500), (41213,-0.393362), (41214,-0.488995), (41215,-0.647332), (41216,-0.375079), (41217,-0.516691), (41218,-0.169662), (41219,-0.319633), (41220,-0.172795), (41221,-0.336706), (41222,-0.295308), (41223,-0.476406), (41224,-0.380664), (41225,-0.496265), (41226,-0.157595), (41227,-0.340083), (41228,-0.320050), (41229,-0.451913), (41230,-0.535461), (41231,-0.714236), (41232,-0.447093), (41233,-0.586852), (41234,-0.257931), (41235,-0.411622), (41236,-0.260608), (41237,-0.387355), (41238,-0.351536), (41239,-0.517763), (41240,-0.464293), (41241,-0.516727), (41242,-0.254229), (41243,-0.288542), (41244,-0.459421), (41245,-0.473295), (41246,-0.660430), (41247,-0.387250), (41248,-0.535832), (41249,-0.570614), (41250,-0.323445), (41251,-0.180327), (41252,-0.357706), (41253,-0.404567), (41254,-0.516448), (41255,-0.220507), (41256,-0.381631), (41257,-0.433132), (41258,-0.232419), (41259,-0.214245), (41260,-0.384192), (41261,-0.431979), (41262,-0.637692), (41263,-0.315741), (41264,-0.487547), (41265,-0.520932), (41266,-0.319286), (41267,-0.176631), (41268,-0.333108), (41269,-0.341410), (41270,-0.430537), (41271,-0.111841), (41272,-0.498704), (41273,-0.524663), (41274,-0.270989), (41275,-0.241207), (41276,-0.406044), (41277,-0.454758), (41278,-0.623314), (41279,-0.332483), (41280,-0.481528), (41281,-0.558112), (41282,-0.312804), (41283,-0.182227), (41284,-0.333126), (41285,-0.389279), (41286,-0.451925), (41287,-0.172709), (41288,-0.414652), (41289,-0.471262), (41290,-0.235709), (41291,-0.226359), (41292,-0.384233), (41293,-0.444562), (41294,-0.649812), (41295,-0.334360), (41296,-0.510349), (41297,-0.574855), (41298,-0.323973), (41299,-0.170635), (41300,-0.349404), (41301,-0.418557), (41302,-0.498861), (41303,-0.185732), (41304,-0.448583), (41305,-0.493114), (41306,-0.290541), (41307,-0.250534), (41308,-0.393542), (41309,-0.460371), (41310,-0.611739), (41311,-0.345066), (41312,-0.515012), (41313,-0.568836), (41314,-0.338392), (41315,-0.184585), (41316,-0.298796), (41317,-0.360979), (41318,-0.393438), (41319,-0.146739), (41320,-0.488549), (41321,-0.172634), (41322,-0.296131), (41323,-0.310012), (41324,-0.460916), (41325,-0.548647), (41326,-0.675864), (41327,-0.410117), (41328,-0.599574), (41329,-0.259508), (41330,-0.403906), (41331,-0.259855), (41332,-0.416796), (41333,-0.400019), (41334,-0.518407), (41335,-0.268452), (41336,-0.456056), (41337,-0.489905), (41338,-0.248773), (41339,-0.204589), (41340,-0.365712), (41341,-0.424182), (41342,-0.609927), (41343,-0.358575), (41344,-0.490438), (41345,-0.645519), (41346,-0.328214), (41347,-0.476332), (41348,-0.345749), (41349,-0.502697), (41350,-0.455720), (41351,-0.632635), (41352,-0.463969), (41353,-0.592576), (41354,-0.297105), (41355,-0.424785), (41356,-0.416361), (41357,-0.564016), (41358,-0.642924), (41359,-0.763635), (41360,-0.521576), (41361,-0.666444), (41362,-0.325444), (41363,-0.464277), (41364,-0.316975), (41365,-0.471593), (41366,-0.431592), (41367,-0.588070), (41368,-0.878785), (41369,-0.581917), (41370,-0.320347), (41371,-0.363025), (41372,-0.489308), (41373,-0.494360), (41374,-0.683354), (41375,-0.742287), (41376,-0.942897), (41377,-0.634878), (41378,-0.394678), (41379,-0.456398), (41380,-0.620308), (41381,-0.457678), (41382,-0.529617), (41383,-0.537455), (41384,-0.910856), (41385,-0.241462), (41386,-0.357064), (41387,-0.436435), (41388,-0.625429), (41389,-0.629084), (41390,-0.753515), (41391,-0.852398), (41392,-0.998656), (41393,-0.313934), (41394,-0.495959), (41395,-0.545600), (41396,-0.717406), (41397,-0.464665), (41398,-0.596528), (41399,-0.618298), (41400,-0.767812), (41401,-0.489060), (41402,-0.259543), (41403,-0.314293), (41404,-0.486099), (41405,-0.481865), (41406,-0.675036), (41407,-0.720500), (41408,-0.855613), (41409,-0.581963), (41410,-0.329222), (41411,-0.369113), (41412,-0.527914), (41413,-0.330914), (41414,-0.436760), (41415,-0.509631), (41416,-0.715344), (41417,-0.403148), (41418,-0.208001), (41419,-0.225595), (41420,-0.400651), (41421,-0.358327), (41422,-0.551034), (41423,-0.641558), (41424,-0.807785), (41425,-0.509064), (41426,-0.295339), (41427,-0.315719), (41428,-0.496347), (41429,-0.310956), (41430,-0.394047), (41431,-0.433469), (41432,-0.850069), (41433,-0.587108), (41434,-0.362231), (41435,-0.395623), (41436,-0.538625), (41437,-0.506057), (41438,-0.692728), (41439,-0.744692), (41440,-0.869122), (41441,-0.588974), (41442,-0.349237), (41443,-0.433255), (41444,-0.588336), (41445,-0.430816), (41446,-0.508334), (41447,-0.553798), (41448,-0.732104), (41449,-0.486795), (41450,-0.191787), (41451,-0.233995), (41452,-0.384900), (41453,-0.376482), (41454,-0.567330), (41455,-0.627197), (41456,-0.786924), (41457,-0.507708), (41458,-0.265185), (41459,-0.335734), (41460,-0.487565), (41461,-0.298925), (41462,-0.395015), (41463,-0.438619), (41464,-0.641082), (41465,-0.365116), (41466,-0.137459), (41467,-0.197319), (41468,-0.365412), (41469,-0.345379), (41470,-0.489321), (41471,-0.584484), (41472,-0.721914), (41473,-0.429692), (41474,-0.221077), (41475,-0.250749), (41476,-0.439274), (41477,-0.271535), (41478,-0.338370), (41479,-0.420991), (41480,-0.761412), (41481,-0.450142), (41482,-0.222479), (41483,-0.299996), (41484,-0.443005), (41485,-0.394638), (41486,-0.550652), (41487,-0.594720), (41488,-0.758631), (41489,-0.499853), (41490,-0.272659), (41491,-0.319050), (41492,-0.471345), (41493,-0.314757), (41494,-0.383446), (41495,-0.425654), (41496,-0.244446), (41497,-0.378626), (41498,-0.435242), (41499,-0.211298), (41500,-0.172687), (41501,-0.333811), (41502,-0.380202), (41503,-0.553868), (41504,-0.291371), (41505,-0.468286), (41506,-0.499349), (41507,-0.285160), (41508,-0.129963), (41509,-0.281794), (41510,-0.345374), (41511,-0.389448), (41512,-0.376848), (41513,-0.562586), (41514,-0.204874), (41515,-0.351132), (41516,-0.382195), (41517,-0.527527), (41518,-0.587850), (41519,-0.708561), (41520,-0.448393), (41521,-0.631345), (41522,-0.288028), (41523,-0.463084), (41524,-0.283266), (41525,-0.445786), (41526,-0.362116), (41527,-0.522313), (41528,-0.323916), (41529,-0.493399), (41530,-0.195599), (41531,-0.371124), (41532,-0.394291), (41533,-0.521044), (41534,-0.618067), (41535,-0.753637), (41536,-0.466989), (41537,-0.625326), (41538,-0.294551), (41539,-0.423158), (41540,-0.270747), (41541,-0.414683), (41542,-0.389540), (41543,-0.558560), (41544,-0.394077), (41545,-0.543585), (41546,-0.200732), (41547,-0.338631), (41548,-0.320458), (41549,-0.484368), (41550,-0.566989), (41551,-0.756447), (41552,-0.450287), (41553,-0.605375), (41554,-0.254156), (41555,-0.380446), (41556,-0.255906), (41557,-0.373830), (41558,-0.351474), (41559,-0.535823), (41560,-0.206438), (41561,-0.361989), (41562,-0.418599), (41563,-0.190942), (41564,-0.158837), (41565,-0.329710), (41566,-0.390966), (41567,-0.558126), (41568,-0.268228), (41569,-0.390798), (41570,-0.439976), (41571,-0.199776), (41572,-0.075699), (41573,-0.234500), (41574,-0.276245), (41575,-0.351903), (41576,-0.389008), (41577,-0.168777), (41578,-0.231893), (41579,-0.386048), (41580,-0.352083), (41581,-0.542004), (41582,-0.579109), (41583,-0.743019), (41584,-0.449401), (41585,-0.211988), (41586,-0.311798), (41587,-0.468275), (41588,-0.303322), (41589,-0.356219), (41590,-0.418402), (41591,-0.609720), (41592,-0.312383), (41593,-0.460037), (41594,-0.125080), (41595,-0.312678), (41596,-0.301938), (41597,-0.439373), (41598,-0.523391), (41599,-0.699837), (41600,-0.669591), (41601,-0.818636), (41602,-0.487398), (41603,-0.624828), (41604,-0.501684), (41605,-0.637724), (41606,-0.600972), (41607,-0.756980), (41608,-0.471265), (41609,-0.607768), (41610,-0.289529), (41611,-0.387485), (41612,-0.358160), (41613,-0.510461), (41614,-0.583326), (41615,-0.741200), (41616,-0.462911), (41617,-0.615206), (41618,-0.289077), (41619,-0.407465), (41620,-0.315905), (41621,-0.465877), (41622,-0.413797), (41623,-0.590712), (41624,-0.852167), (41625,-0.574341), (41626,-0.311850), (41627,-0.367527), (41628,-0.503567), (41629,-0.459389), (41630,-0.649310), (41631,-0.717529), (41632,-0.861465), (41633,-0.588755), (41634,-0.350872), (41635,-0.390764), (41636,-0.534236), (41637,-0.412945), (41638,-0.482561), (41639,-0.551720), (41640,-0.764865), (41641,-0.507941), (41642,-0.263559), (41643,-0.291371), (41644,-0.472470), (41645,-0.436182), (41646,-0.629816), (41647,-0.681786), (41648,-0.834081), (41649,-0.522818), (41650,-0.312343), (41651,-0.357807), (41652,-0.555624), (41653,-0.409713), (41654,-0.483981), (41655,-0.553133), (41656,-0.949752), (41657,-0.656598), (41658,-0.414539), (41659,-0.451644), (41660,-0.605798), (41661,-0.569973), (41662,-0.752931), (41663,-0.818364), (41664,-0.990170), (41665,-0.679834), (41666,-0.444281), (41667,-0.485562), (41668,-0.657368), (41669,-0.515640), (41670,-0.562964), (41671,-0.599136), (41672,-0.756077), (41673,-0.458283), (41674,-0.251990), (41675,-0.290022), (41676,-0.439994), (41677,-0.433899), (41678,-0.595950), (41679,-0.666035), (41680,-0.811361), (41681,-0.529822), (41682,-0.260825), (41683,-0.304429), (41684,-0.459047), (41685,-0.301063), (41686,-0.402269), (41687,-0.443551), (41688,-0.865254), (41689,-0.528437), (41690,-0.307286), (41691,-0.348104), (41692,-0.528733), (41693,-0.534254), (41694,-0.696767), (41695,-0.758024), (41696,-0.936336), (41697,-0.679875), (41698,-0.441998), (41699,-0.499535), (41700,-0.635111), (41701,-0.494316), (41702,-0.587156), (41703,-0.588958), (41704,-0.740789), (41705,-0.442525), (41706,-0.235769), (41707,-0.291916), (41708,-0.412164), (41709,-0.435337), (41710,-0.609929), (41711,-0.671649), (41712,-0.848564), (41713,-0.540545), (41714,-0.280371), (41715,-0.350919), (41716,-0.484636), (41717,-0.300178), (41718,-0.406023), (41719,-0.450561), (41720,-0.504384), (41721,-0.208444), (41722,-0.349129), (41723,-0.025318), (41724,-0.193874), (41725,-0.194279), (41726,-0.347970), (41727,-0.425488), (41728,-0.639097), (41729,-0.392855), (41730,-0.519145), (41731,-0.178615), (41732,-0.331373), (41733,-0.181749), (41734,-0.325684), (41735,-0.280574), (41736,-0.549924), (41737,-0.262812), (41738,-0.466666), (41739,-0.123812), (41740,-0.268211), (41741,-0.278842), (41742,-0.389334), (41743,-0.475674), (41744,-0.615890), (41745,-0.336211), (41746,-0.480146), (41747,-0.177706), (41748,-0.307703), (41749,-0.151115), (41750,-0.299697), (41751,-0.293133), (41752,-0.234553), (41753,-0.379416), (41754,-0.441141), (41755,-0.161919), (41756,-0.169764), (41757,-0.309516), (41758,-0.391210), (41759,-0.567663), (41760,-0.294946), (41761,-0.429596), (41762,-0.492706), (41763,-0.257152), (41764,-0.100559), (41765,-0.301632), (41766,-0.312256), (41767,-0.368866), (41768,-0.339548), (41769,-0.519713), (41770,-0.149922), (41771,-0.297571), (41772,-0.288690), (41773,-0.425199), (41774,-0.514320), (41775,-0.666621), (41776,-0.421312), (41777,-0.616806), (41778,-0.269770), (41779,-0.400700), (41780,-0.271977), (41781,-0.407089), (41782,-0.383344), (41783,-0.496622), (41784,-0.191858), (41785,-0.372957), (41786,-0.414238), (41787,-0.185648), (41788,-0.183736), (41789,-0.349506), (41790,-0.394038), (41791,-0.576063), (41792,-0.290804), (41793,-0.441246), (41794,-0.474631), (41795,-0.239541), (41796,-0.104782), (41797,-0.239432), (41798,-0.275604), (41799,-0.352652), (41800,-0.157042), (41801,-0.329311), (41802,-0.390104), (41803,-0.128540), (41804,-0.105721), (41805,-0.248729), (41806,-0.315559), (41807,-0.528241), (41808,-0.223477), (41809,-0.386455), (41810,-0.420773), (41811,-0.208908), (41812,-0.048131), (41813,-0.202756), (41814,-0.245433), (41815,-0.304830), (41816,-0.175180), (41817,-0.352559), (41818,-0.357611), (41819,-0.146672), (41820,-0.141505), (41821,-0.297982), (41822,-0.343916), (41823,-0.529655), (41824,-0.236037), (41825,-0.377186), (41826,-0.405462), (41827,-0.166659), (41828,-0.047228), (41829,-0.201846), (41830,-0.246377), (41831,-0.315066), (41832,-0.236049), (41833,-0.412501), (41834,-0.079397), (41835,-0.205687), (41836,-0.211665), (41837,-0.354211), (41838,-0.440081), (41839,-0.605388), (41840,-0.363329), (41841,-0.504014), (41842,-0.155588), (41843,-0.328321), (41844,-0.114596), (41845,-0.284542), (41846,-0.265906), (41847,-0.416811), (41848,-0.435337), (41849,-0.554188), (41850,-0.210872), (41851,-0.383605), (41852,-0.388193), (41853,-0.555359), (41854,-0.630084), (41855,-0.820005), (41856,-0.524991), (41857,-0.681938), (41858,-0.706032), (41859,-0.426352), (41860,-0.303666), (41861,-0.491733), (41862,-0.550197), (41863,-0.609136), (41864,-0.893809), (41865,-0.581613), (41866,-0.379503), (41867,-0.394774), (41868,-0.533600), (41869,-0.542371), (41870,-0.686769), (41871,-0.728521), (41872,-0.852018), (41873,-0.574655), (41874,-0.340962), (41875,-0.370165), (41876,-0.546617), (41877,-0.433223), (41878,-0.524209), (41879,-0.561308), (41880,-0.655545), (41881,-0.389798), (41882,-0.580652), (41883,-0.230829), (41884,-0.364546), (41885,-0.347306), (41886,-0.512606), (41887,-0.562253), (41888,-0.710835), (41889,-0.485031), (41890,-0.587627), (41891,-0.284253), (41892,-0.428195), (41893,-0.274388), (41894,-0.460596), (41895,-0.424308), (41896,-0.840901), (41897,-0.549607), (41898,-0.320553), (41899,-0.395278), (41900,-0.580090), (41901,-0.552631), (41902,-0.728619), (41903,-0.755036), (41904,-0.883179), (41905,-0.610000), (41906,-0.385592), (41907,-0.429197), (41908,-0.553164), (41909,-0.407716), (41910,-0.490807), (41911,-0.529765), (41912,-0.751740), (41913,-0.507821), (41914,-0.646183), (41915,-0.268960), (41916,-0.433333), (41917,-0.409124), (41918,-0.547017), (41919,-0.658905), (41920,-0.774506), (41921,-0.516655), (41922,-0.636903), (41923,-0.337249), (41924,-0.477471), (41925,-0.368253), (41926,-0.519621), (41927,-0.502381), (41928,-0.829790), (41929,-0.534782), (41930,-0.287613), (41931,-0.352119), (41932,-0.490482), (41933,-0.433762), (41934,-0.631579), (41935,-0.705378), (41936,-0.864642), (41937,-0.588212), (41938,-0.327105), (41939,-0.394404), (41940,-0.558777), (41941,-0.408220), (41942,-0.447185), (41943,-0.513087), (41944,-0.707185), (41945,-0.435865), (41946,-0.626249), (41947,-0.258312), (41948,-0.444056), (41949,-0.412415), (41950,-0.560063), (41951,-0.660342), (41952,-0.756895), (41953,-0.471643), (41954,-0.628121), (41955,-0.282011), (41956,-0.453818), (41957,-0.289334), (41958,-0.420728), (41959,-0.411847), (41960,-0.537667), (41961,-0.300718), (41962,-0.500395), (41963,-0.136640), (41964,-0.264314), (41965,-0.251256), (41966,-0.403551), (41967,-0.491751), (41968,-0.670984), (41969,-0.382476), (41970,-0.536167), (41971,-0.175198), (41972,-0.355370), (41973,-0.193204), (41974,-0.353858), (41975,-0.312466), (41976,-0.507027), (41977,-0.244067), (41978,-0.404727), (41979,-0.073953), (41980,-0.248545), (41981,-0.211330), (41982,-0.391959), (41983,-0.449033), (41984,-0.583682), (41985,-0.362524), (41986,-0.499960), (41987,-0.179398), (41988,-0.370716), (41989,-0.204373), (41990,-0.386861), (41991,-0.371012), (41992,-0.701676), (41993,-0.382048), (41994,-0.585438), (41995,-0.199385), (41996,-0.334498), (41997,-0.344659), (41998,-0.442145), (41999,-0.470884), (42000,-0.683103), (42001,-0.396918), (42002,-0.551073), (42003,-0.189178), (42004,-0.359587), (42005,-0.244803), (42006,-0.416146), (42007,-0.377535), (42008,-0.384909), (42009,-0.535351), (42010,-0.611935), (42011,-0.320641), (42012,-0.333588), (42013,-0.469164), (42014,-0.525774), (42015,-0.718945), (42016,-0.439729), (42017,-0.585061), (42018,-0.645384), (42019,-0.407508), (42020,-0.269499), (42021,-0.406002), (42022,-0.459362), (42023,-0.542916), (42024,-0.292492), (42025,-0.453152), (42026,-0.495830), (42027,-0.252381), (42028,-0.267651), (42029,-0.374424), (42030,-0.420821), (42031,-0.638613), (42032,-0.307832), (42033,-0.479175), (42034,-0.517206), (42035,-0.283976), (42036,-0.117164), (42037,-0.247630), (42038,-0.304240), (42039,-0.385935), (42040,-0.246066), (42041,-0.398824), (42042,-0.458690), (42043,-0.240319), (42044,-0.210074), (42045,-0.357722), (42046,-0.418052), (42047,-0.596364), (42048,-0.310179), (42049,-0.457827), (42050,-0.493999), (42051,-0.239404), (42052,-0.109748), (42053,-0.282487), (42054,-0.331665), (42055,-0.426365), (42056,-0.249803), (42057,-0.373763), (42058,-0.387644), (42059,-0.162303), (42060,-0.183153), (42061,-0.344740), (42062,-0.378589), (42063,-0.587089), (42064,-0.271643), (42065,-0.426261), (42066,-0.494023), (42067,-0.275651), (42068,-0.099553), (42069,-0.278328), (42070,-0.325183), (42071,-0.396195), (42072,-0.278617), (42073,-0.458789), (42074,-0.502394), (42075,-0.268694), (42076,-0.271429), (42077,-0.421400), (42078,-0.452932), (42079,-0.657249), (42080,-0.366888), (42081,-0.554486), (42082,-0.588798), (42083,-0.323984), (42084,-0.165067), (42085,-0.331764), (42086,-0.402312), (42087,-0.484470), (42088,-0.738029), (42089,-0.443478), (42090,-0.188883), (42091,-0.238060), (42092,-0.398251), (42093,-0.361500), (42094,-0.540738), (42095,-0.599672), (42096,-0.762655), (42097,-0.491798), (42098,-0.258099), (42099,-0.253401), (42100,-0.420561), (42101,-0.259321), (42102,-0.345661), (42103,-0.411101), (42104,-0.273549), (42105,-0.450001), (42106,-0.525196), (42107,-0.295215), (42108,-0.266360), (42109,-0.414942), (42110,-0.434852), (42111,-0.612237), (42112,-0.782647), (42113,-0.523869), (42114,-0.678024), (42115,-0.327738), (42116,-0.499081), (42117,-0.373607), (42118,-0.491068), (42119,-0.464536), (42120,-0.704626), (42121,-0.415185), (42122,-0.572595), (42123,-0.211157), (42124,-0.380640), (42125,-0.362004), (42126,-0.531956), (42127,-0.611328), (42128,-0.777561), (42129,-0.457932), (42130,-0.622769), (42131,-0.278519), (42132,-0.431747), (42133,-0.258898), (42134,-0.421412), (42135,-0.432506), (42136,-0.672596), (42137,-0.407775), (42138,-0.569363), (42139,-0.231619), (42140,-0.398315), (42141,-0.398257), (42142,-0.577033), (42143,-0.636893), (42144,-0.775718), (42145,-0.519264), (42146,-0.661339), (42147,-0.338461), (42148,-0.494938), (42149,-0.327662), (42150,-0.428868), (42151,-0.417664), (42152,-0.735787), (42153,-0.883436), (42154,-0.234017), (42155,-0.336150), (42156,-0.400192), (42157,-0.554347), (42158,-0.577513), (42159,-0.738637), (42160,-0.816618), (42161,-0.960090), (42162,-0.256790), (42163,-0.418840), (42164,-0.492639), (42165,-0.608240), (42166,-0.407984), (42167,-0.564462), (42168,-0.741377), (42169,-0.475167), (42170,-0.625145), (42171,-0.301333), (42172,-0.468030), (42173,-0.452643), (42174,-0.581713), (42175,-0.661554), (42176,-0.801307), (42177,-0.556461), (42178,-0.704116), (42179,-0.390987), (42180,-0.532142), (42181,-0.326777), (42182,-0.549678), (42183,-0.534291), (42184,-0.597871), (42185,-0.745056), (42186,-0.467700), (42187,-0.246542), (42188,-0.295719), (42189,-0.433155), (42190,-0.428451), (42191,-0.591898), (42192,-0.662910), (42193,-0.837966), (42194,-0.522520), (42195,-0.301362), (42196,-0.330102), (42197,-0.510737), (42198,-0.342071), (42199,-0.428405), (42200,-0.760929), (42201,-0.497036), (42202,-0.638654), (42203,-0.288832), (42204,-0.440663), (42205,-0.414131), (42206,-0.555743), (42207,-0.630938), (42208,-0.795775), (42209,-0.526315), (42210,-0.692078), (42211,-0.331110), (42212,-0.473192), (42213,-0.350969), (42214,-0.519988), (42215,-0.483700), (42216,-0.524518), (42217,-0.659631), (42218,-0.363227), (42219,-0.143466), (42220,-0.182887), (42221,-0.326359), (42222,-0.342100), (42223,-0.493931), (42224,-0.537999), (42225,-0.728390), (42226,-0.447777), (42227,-0.214078), (42228,-0.256756), (42229,-0.468975), (42230,-0.304948), (42231,-0.364345), (42232,-0.687577), (42233,-0.442731), (42234,-0.566698), (42235,-0.206193), (42236,-0.357561), (42237,-0.318487), (42238,-0.438271), (42239,-0.577560), (42240,-0.682016), (42241,-0.391185), (42242,-0.585289), (42243,-0.208992), (42244,-0.383115), (42245,-0.249752), (42246,-0.385791), (42247,-0.356472), (42248,-0.572405), (42249,-0.707981), (42250,-0.463598), (42251,-0.238264), (42252,-0.263754), (42253,-0.442529), (42254,-0.440148), (42255,-0.593839), (42256,-0.639767), (42257,-0.773947), (42258,-0.520278), (42259,-0.292151), (42260,-0.348768), (42261,-0.506172), (42262,-0.317995), (42263,-0.399689), (42264,-0.666253), (42265,-0.408865), (42266,-0.559770), (42267,-0.273585), (42268,-0.419843), (42269,-0.382165), (42270,-0.497766), (42271,-0.592466), (42272,-0.745694), (42273,-0.453003), (42274,-0.624809), (42275,-0.268017), (42276,-0.389661), (42277,-0.257689), (42278,-0.416489), (42279,-0.383914), (42280,-0.583128), (42281,-0.299729), (42282,-0.476181), (42283,-0.151906), (42284,-0.262398), (42285,-0.256304), (42286,-0.405812), (42287,-0.494476), (42288,-0.662105), (42289,-0.389389), (42290,-0.542147), (42291,-0.205337), (42292,-0.334407), (42293,-0.223335), (42294,-0.313853), (42295,-0.283144), (42296,-0.626814), (42297,-0.379176), (42298,-0.534726), (42299,-0.215098), (42300,-0.343241), (42301,-0.337147), (42302,-0.495947), (42303,-0.588324), (42304,-0.711822), (42305,-0.455830), (42306,-0.588157), (42307,-0.270381), (42308,-0.414786), (42309,-0.262376), (42310,-0.411884), (42311,-0.399753), (42312,-0.674207), (42313,-0.390345), (42314,-0.529640), (42315,-0.204432), (42316,-0.358593), (42317,-0.370608), (42318,-0.479709), (42319,-0.548398), (42320,-0.686761), (42321,-0.426123), (42322,-0.581204), (42323,-0.258789), (42324,-0.405517), (42325,-0.257283), (42326,-0.412371), (42327,-0.393265), (42328,-0.618489), (42329,-0.355065), (42330,-0.511079), (42331,-0.170086), (42332,-0.316808), (42333,-0.313963), (42334,-0.480660), (42335,-0.535880), (42336,-0.733233), (42337,-0.434037), (42338,-0.574722), (42339,-0.288537), (42340,-0.432009), (42341,-0.278672), (42342,-0.441655), (42343,-0.379356), (42344,-0.731849), (42345,-0.441018), (42346,-0.225902), (42347,-0.282976), (42348,-0.437130), (42349,-0.441255), (42350,-0.576368), (42351,-0.618576), (42352,-0.764835), (42353,-0.502807), (42354,-0.261211), (42355,-0.311785), (42356,-0.461757), (42357,-0.322351), (42358,-0.377108), (42359,-0.420249), (42360,-0.607847), (42361,-0.336064), (42362,-0.506474), (42363,-0.151078), (42364,-0.303843), (42365,-0.287993), (42366,-0.456549), (42367,-0.524305), (42368,-0.759749), (42369,-0.453589), (42370,-0.620285), (42371,-0.293224), (42372,-0.437623), (42373,-0.293114), (42374,-0.477456), (42375,-0.401688), (42376,-0.821068), (42377,-0.556718), (42378,-0.302580), (42379,-0.344794), (42380,-0.502199), (42381,-0.469167), (42382,-0.604743), (42383,-0.651134), (42384,-0.833622), (42385,-0.542791), (42386,-0.337895), (42387,-0.389395), (42388,-0.534264), (42389,-0.400895), (42390,-0.520216), (42391,-0.531767), (42392,-0.534965), (42393,-0.705375), (42394,-0.410367), (42395,-0.174807), (42396,-0.231424), (42397,-0.399047), (42398,-0.407818), (42399,-0.539674), (42400,-0.567950), (42401,-0.743939), (42402,-0.468900), (42403,-0.211982), (42404,-0.275555), (42405,-0.430642), (42406,-0.282878), (42407,-0.341811), (42408,-0.651568), (42409,-0.829417), (42410,-0.158164), (42411,-0.329043), (42412,-0.398659), (42413,-0.540734), (42414,-0.569943), (42415,-0.728281), (42416,-0.777922), (42417,-0.960880), (42418,-0.309138), (42419,-0.461433), (42420,-0.471131), (42421,-0.606243), (42422,-0.373940), (42423,-0.518339), (42424,-0.565193), (42425,-0.735146), (42426,-0.465679), (42427,-0.237559), (42428,-0.274657), (42429,-0.434391), (42430,-0.438979), (42431,-0.597310), (42432,-0.669718), (42433,-0.834555), (42434,-0.522359), (42435,-0.309561), (42436,-0.356421), (42437,-0.504540), (42438,-0.349806), (42439,-0.394801), (42440,-0.628384), (42441,-0.796477), (42442,-0.134053), (42443,-0.285421), (42444,-0.345281), (42445,-0.505015), (42446,-0.523072), (42447,-0.653538), (42448,-0.697606), (42449,-0.874522), (42450,-0.199556), (42451,-0.338382), (42452,-0.393138), (42453,-0.556579), (42454,-0.300124), (42455,-0.453352), (42456,-0.554088), (42457,-0.683158), (42458,-0.437849), (42459,-0.200436), (42460,-0.199452), (42461,-0.365221), (42462,-0.350298), (42463,-0.520714), (42464,-0.559673), (42465,-0.778855), (42466,-0.493133), (42467,-0.222276), (42468,-0.293288), (42469,-0.454875), (42470,-0.270881), (42471,-0.370690), (42472,-0.383637), (42473,-0.546158), (42474,-0.267868), (42475,-0.042991), (42476,-0.061055), (42477,-0.259335), (42478,-0.265783), (42479,-0.454308), (42480,-0.479797), (42481,-0.657183), (42482,-0.384466), (42483,-0.139621), (42484,-0.176256), (42485,-0.342026), (42486,-0.210980), (42487,-0.288028), (42488,-0.443116), (42489,-0.610739), (42490,-0.312945), (42491,-0.086214), (42492,-0.133532), (42493,-0.290942), (42494,-0.234216), (42495,-0.419955), (42496,-0.523947), (42497,-0.675778), (42498,-0.373801), (42499,-0.099695), (42500,-0.206004), (42501,-0.383852), (42502,-0.216113), (42503,-0.265290), (42504,-0.484472), (42505,-0.666034), (42506,-0.379386), (42507,-0.127571), (42508,-0.166999), (42509,-0.334622), (42510,-0.311809), (42511,-0.485469), (42512,-0.556481), (42513,-0.669759), (42514,-0.375678), (42515,-0.137338), (42516,-0.221819), (42517,-0.377833), (42518,-0.187796), (42519,-0.284819), (42520,-0.529549), (42521,-0.254516), (42522,-0.413780), (42523,-0.102973), (42524,-0.242269), (42525,-0.246387), (42526,-0.444674), (42527,-0.518003), (42528,-0.691206), (42529,-0.406880), (42530,-0.537810), (42531,-0.211212), (42532,-0.334709), (42533,-0.215279), (42534,-0.353178), (42535,-0.321999), (42536,-0.522140), (42537,-0.272184), (42538,-0.424949), (42539,-0.070017), (42540,-0.228354), (42541,-0.227833), (42542,-0.388487), (42543,-0.472504), (42544,-0.576033), (42545,-0.313536), (42546,-0.470477), (42547,-0.135519), (42548,-0.304076), (42549,-0.141909), (42550,-0.296990), (42551,-0.255599), (42552,-0.622024), (42553,-0.351631), (42554,-0.497889), (42555,-0.151323), (42556,-0.318946), (42557,-0.294274), (42558,-0.413125), (42559,-0.472991), (42560,-0.647120), (42561,-0.371618), (42562,-0.546673), (42563,-0.205217), (42564,-0.377486), (42565,-0.227398), (42566,-0.338353), (42567,-0.313681), (42568,-0.548191), (42569,-0.285231), (42570,-0.390150), (42571,-0.070984), (42572,-0.220962), (42573,-0.236233), (42574,-0.394100), (42575,-0.487410), (42576,-0.637851), (42577,-0.353056), (42578,-0.498852), (42579,-0.140670), (42580,-0.312012), (42581,-0.162851), (42582,-0.302610), (42583,-0.290010), (42584,-0.556111), (42585,-0.255060), (42586,-0.415714), (42587,-0.089586), (42588,-0.250247), (42589,-0.231610), (42590,-0.399697), (42591,-0.456307), (42592,-0.604425), (42593,-0.310344), (42594,-0.458926), (42595,-0.151839), (42596,-0.302744), (42597,-0.159619), (42598,-0.325389), (42599,-0.295607), (42600,-0.642063), (42601,-0.355408), (42602,-0.150049), (42603,-0.187611), (42604,-0.344558), (42605,-0.343104), (42606,-0.540921), (42607,-0.534363), (42608,-0.741009), (42609,-0.445532), (42610,-0.211369), (42611,-0.235005), (42612,-0.417957), (42613,-0.252077), (42614,-0.327266), (42615,-0.381089), (42616,-0.553829), (42617,-0.257424), (42618,-0.398573), (42619,-0.060360), (42620,-0.192223), (42621,-0.240010), (42622,-0.428998), (42623,-0.488865), (42624,-0.781440), (42625,-0.504077), (42626,-0.678206), (42627,-0.352078), (42628,-0.469069), (42629,-0.317122), (42630,-0.479179), (42631,-0.437781), (42632,-0.678797), (42633,-0.391679), (42634,-0.549090), (42635,-0.185335), (42636,-0.378506), (42637,-0.366369), (42638,-0.493123), (42639,-0.578067), (42640,-0.733618), (42641,-0.460438), (42642,-0.580685), (42643,-0.223430), (42644,-0.401742), (42645,-0.248862), (42646,-0.415095), (42647,-0.388563), (42648,-0.565942), (42649,-0.744254), (42650,-0.482683), (42651,-0.198358), (42652,-0.262401), (42653,-0.427244), (42654,-0.399778), (42655,-0.589236), (42656,-0.651419), (42657,-0.812543), (42658,-0.511962), (42659,-0.242959), (42660,-0.314434), (42661,-0.479741), (42662,-0.323147), (42663,-0.365825), (42664,-0.749439), (42665,-0.867826), (42666,-0.169172), (42667,-0.317291), (42668,-0.393875), (42669,-0.575437), (42670,-0.553081), (42671,-0.709096), (42672,-0.783821), (42673,-0.922183), (42674,-0.238394), (42675,-0.390689), (42676,-0.451482), (42677,-0.603313), (42678,-0.370547), (42679,-0.499153), (42680,-0.606859), (42681,-0.793993), (42682,-0.491090), (42683,-0.251354), (42684,-0.294025), (42685,-0.459795), (42686,-0.472743), (42687,-0.651518), (42688,-0.703952), (42689,-0.883190), (42690,-0.597005), (42691,-0.373061), (42692,-0.413416), (42693,-0.606123), (42694,-0.426305), (42695,-0.482915), (42696,-0.540922), (42697,-0.696936), (42698,-0.434902), (42699,-0.197952), (42700,-0.290799), (42701,-0.411973), (42702,-0.356180), (42703,-0.536345), (42704,-0.587846), (42705,-0.767548), (42706,-0.497618), (42707,-0.281576), (42708,-0.276409), (42709,-0.429637), (42710,-0.273043), (42711,-0.372389), (42712,-0.605973), (42713,-0.761524), (42714,-0.466509), (42715,-0.234206), (42716,-0.278274), (42717,-0.410137), (42718,-0.420298), (42719,-0.597214), (42720,-0.655220), (42721,-0.791723), (42722,-0.543164), (42723,-0.306678), (42724,-0.309870), (42725,-0.466347), (42726,-0.372928), (42727,-0.424898), (42728,-0.490331), (42729,-0.648668), (42730,-0.369452), (42731,-0.122747), (42732,-0.135694), (42733,-0.300068), (42734,-0.315808), (42735,-0.477858), (42736,-0.514030), (42737,-0.677014), (42738,-0.373640), (42739,-0.167811), (42740,-0.210489), (42741,-0.367900), (42742,-0.222452), (42743,-0.264666), (42744,-0.449941), (42745,-0.592487), (42746,-0.308155), (42747,-0.062383), (42748,-0.139894), (42749,-0.305201), (42750,-0.271699), (42751,-0.474162), (42752,-0.540065), (42753,-0.685860), (42754,-0.411284), (42755,-0.179914), (42756,-0.212366), (42757,-0.407866), (42758,-0.214579), (42759,-0.258647), (42760,-0.491768), (42761,-0.654745), (42762,-0.388071), (42763,-0.183638), (42764,-0.195659), (42765,-0.371642), (42766,-0.379949), (42767,-0.570334), (42768,-0.620908), (42769,-0.747192), (42770,-0.448464), (42771,-0.234276), (42772,-0.266271), (42773,-0.446437), (42774,-0.287057), (42775,-0.355282), (42776,-0.621846), (42777,-0.335198), (42778,-0.479133), (42779,-0.152072), (42780,-0.292757), (42781,-0.297809), (42782,-0.427349), (42783,-0.509970), (42784,-0.645083), (42785,-0.397451), (42786,-0.520015), (42787,-0.167412), (42788,-0.358260), (42789,-0.165900), (42790,-0.320061), (42791,-0.316753), (42792,-0.496918), (42793,-0.244640), (42794,-0.409013), (42795,-0.036430), (42796,-0.175262), (42797,-0.185886), (42798,-0.379057), (42799,-0.454715), (42800,-0.592151), (42801,-0.322685), (42802,-0.501460), (42803,-0.152101), (42804,-0.316938), (42805,-0.147808), (42806,-0.321474), (42807,-0.301905), (42808,-0.619101), (42809,-0.312477), (42810,-0.478241), (42811,-0.151649), (42812,-0.278396), (42813,-0.267193), (42814,-0.405555), (42815,-0.536022), (42816,-0.648837), (42817,-0.386339), (42818,-0.558609), (42819,-0.180458), (42820,-0.314175), (42821,-0.205427), (42822,-0.342393), (42823,-0.312611), (42824,-0.563383), (42825,-0.294843), (42826,-0.470832), (42827,-0.114973), (42828,-0.272847), (42829,-0.261637), (42830,-0.434839), (42831,-0.475194), (42832,-0.624702), (42833,-0.384503), (42834,-0.525652), (42835,-0.172116), (42836,-0.349495), (42837,-0.198481), (42838,-0.348453), (42839,-0.335852), (42840,-0.585698), (42841,-0.299049), (42842,-0.433692), (42843,-0.091302), (42844,-0.238494), (42845,-0.237503), (42846,-0.408846), (42847,-0.485430), (42848,-0.667456), (42849,-0.375234), (42850,-0.495945), (42851,-0.179103), (42852,-0.329081), (42853,-0.198498), (42854,-0.347080), (42855,-0.316828), (42856,-0.648426), (42857,-0.380819), (42858,-0.138760), (42859,-0.186547), (42860,-0.338842), (42861,-0.292798), (42862,-0.507804), (42863,-0.540726), (42864,-0.700459), (42865,-0.417987), (42866,-0.186147), (42867,-0.185163), (42868,-0.372761), (42869,-0.227319), (42870,-0.296935), (42871,-0.341936), (42872,-0.552758), (42873,-0.315345), (42874,-0.431410), (42875,-0.080197), (42876,-0.253394), (42877,-0.213856), (42878,-0.388448), (42879,-0.447381), (42880,-0.720451), (42881,-0.456094), (42882,-0.581451), (42883,-0.230702), (42884,-0.407618), (42885,-0.241738), (42886,-0.383351), (42887,-0.367501), (42888,-0.618273), (42889,-0.326515), (42890,-0.511790), (42891,-0.128987), (42892,-0.284538), (42893,-0.269151), (42894,-0.431671), (42895,-0.501750), (42896,-0.658228), (42897,-0.395730), (42898,-0.554068), (42899,-0.253950), (42900,-0.410428), (42901,-0.231536), (42902,-0.365259), (42903,-0.309460), (42904,-0.555586), (42905,-0.702771), (42906,-0.427738), (42907,-0.201007), (42908,-0.274806), (42909,-0.422454), (42910,-0.422396), (42911,-0.611854), (42912,-0.672183), (42913,-0.818442), (42914,-0.521574), (42915,-0.300880), (42916,-0.350064), (42917,-0.518150), (42918,-0.393610), (42919,-0.440465), (42920,-0.522159), (42921,-0.703258), (42922,-0.419396), (42923,-0.169440), (42924,-0.215831), (42925,-0.376955), (42926,-0.362032), (42927,-0.558922), (42928,-0.585345), (42929,-0.718135), (42930,-0.454704), (42931,-0.221938), (42932,-0.295273), (42933,-0.460109), (42934,-0.284474), (42935,-0.354090), (42936,-0.591393), (42937,-0.727432), (42938,-0.488160), (42939,-0.205224), (42940,-0.253475), (42941,-0.444329), (42942,-0.449844), (42943,-0.640229), (42944,-0.676870), (42945,-0.844494), (42946,-0.554132), (42947,-0.309286), (42948,-0.356141), (42949,-0.546525), (42950,-0.412693), (42951,-0.483705), (42952,-0.591410), (42953,-0.710268), (42954,-0.441264), (42955,-0.206175), (42956,-0.226555), (42957,-0.359344), (42958,-0.378798), (42959,-0.556640), (42960,-0.581203), (42961,-0.741863), (42962,-0.474720), (42963,-0.223838), (42964,-0.284161), (42965,-0.431816), (42966,-0.292411), (42967,-0.355990), (42968,-0.656461), (42969,-0.812475), (42970,-0.495170), (42971,-0.241495), (42972,-0.268844), (42973,-0.424395), (42974,-0.424337), (42975,-0.601253), (42976,-0.697813), (42977,-0.824560), (42978,-0.557423), (42979,-0.334868), (42980,-0.353858), (42981,-0.537743), (42982,-0.396015), (42983,-0.471203), (42984,-0.565903), (42985,-0.738179), (42986,-0.440842), (42987,-0.193210), (42988,-0.257253), (42989,-0.397012), (42990,-0.394167), (42991,-0.552035), (42992,-0.563592), (42993,-0.699168), (42994,-0.410660), (42995,-0.235951), (42996,-0.308360), (42997,-0.432320), (42998,-0.280843), (42999,-0.354635), (43000,-0.451194), (43001,-0.576088), (43002,-0.308018), (43003,-0.080361), (43004,-0.128142), (43005,-0.309240), (43006,-0.241832), (43007,-0.463806), (43008,-0.906411), (43009,-1.064748), (43010,-0.390709), (43011,-0.489122), (43012,-0.550848), (43013,-0.704069), (43014,-0.455510), (43015,-0.618024), (43016,-0.867869), (43017,-0.998336), (43018,-0.328010), (43019,-0.464049), (43020,-0.549000), (43021,-0.679930), (43022,-0.683585), (43023,-0.856324), (43024,-0.898069), (43025,-1.049900), (43026,-0.390263), (43027,-0.556959), (43028,-0.598710), (43029,-0.790955), (43030,-0.521951), (43031,-0.690508), (43032,-0.783811), (43033,-0.520387), (43034,-0.679188), (43035,-0.340981), (43036,-0.488636), (43037,-0.463030), (43038,-0.608825), (43039,-0.674258), (43040,-0.832132), (43041,-0.537124), (43042,-0.710784), (43043,-0.432494), (43044,-0.551352), (43045,-0.394758), (43046,-0.569351), (43047,-0.517271), (43048,-0.933401), (43049,-0.643503), (43050,-0.400511), (43051,-0.457590), (43052,-0.595953), (43053,-0.616333), (43054,-0.756555), (43055,-0.818738), (43056,-1.001690), (43057,-0.738729), (43058,-0.478555), (43059,-0.535635), (43060,-0.651700), (43061,-0.511831), (43062,-0.541040), (43063,-0.626448), (43064,-0.892548), (43065,-0.632838), (43066,-0.383346), (43067,-0.430207), (43068,-0.595043), (43069,-0.534134), (43070,-0.731025), (43071,-0.782062), (43072,-0.983135), (43073,-0.697413), (43074,-0.419124), (43075,-0.495709), (43076,-0.664729), (43077,-0.516031), (43078,-0.579147), (43079,-0.644117), (43080,-0.918577), (43081,-0.631001), (43082,-0.383833), (43083,-0.452522), (43084,-0.621078), (43085,-0.592686), (43086,-0.777961), (43087,-0.812743), (43088,-0.965037), (43089,-0.671420), (43090,-0.424251), (43091,-0.472038), (43092,-0.583927), (43093,-0.454740), (43094,-0.522966), (43095,-0.599081), (43096,-0.690531), (43097,-0.412242), (43098,-0.580335), (43099,-0.217044), (43100,-0.364229), (43101,-0.343733), (43102,-0.520648), (43103,-0.610708), (43104,-0.744888), (43105,-0.451734), (43106,-0.638405), (43107,-0.289515), (43108,-0.449243), (43109,-0.300082), (43110,-0.472351), (43111,-0.417485), (43112,-0.837335), (43113,-0.590629), (43114,-0.299335), (43115,-0.477640), (43116,-0.514282), (43117,-0.708386), (43118,-0.716687), (43119,-0.885707), (43120,-0.926525), (43121,-0.716983), (43122,-0.411286), (43123,-0.559405), (43124,-0.588614), (43125,-0.654046), (43126,-0.462619), (43127,-0.622346), (43128,-0.837352), (43129,-0.536771), (43130,-0.319790), (43131,-0.371297), (43132,-0.537524), (43133,-0.504955), (43134,-0.701382), (43135,-0.742664), (43136,-1.040348), (43137,-0.835916), (43138,-0.560876), (43139,-0.740115), (43140,-0.773500), (43141,-0.829184), (43142,-0.677236), (43143,-0.846719), (43144,-0.927951), (43145,-0.670099), (43146,-0.392737), (43147,-0.559897), (43148,-0.617440), (43149,-0.757662), (43150,-0.765037), (43151,-0.902466), (43152,-0.953973), (43153,-0.730956), (43154,-0.437338), (43155,-0.632369), (43156,-0.647639), (43157,-0.746522), (43158,-0.616409), (43159,-0.776600), (43160,-0.987422), (43161,-0.756979), (43162,-0.448965), (43163,-0.645386), (43164,-0.714075), (43165,-0.870089), (43166,-0.837051), (43167,-0.985632), (43168,-1.059431), (43169,-0.813195), (43170,-0.539082), (43171,-0.685811), (43172,-0.761926), (43173,-0.827365), (43174,-0.659626), (43175,-0.862552), (43176,-0.913126), (43177,-0.687322), (43178,-0.427618), (43179,-0.551578), (43180,-0.586360), (43181,-0.780464), (43182,-0.793875), (43183,-0.957322), (43184,-0.995354), (43185,-0.760264), (43186,-0.472682), (43187,-0.618477), (43188,-0.676014), (43189,-0.725661), (43190,-0.570927), (43191,-0.747380), (43192,-1.078044), (43193,-0.836912), (43194,-0.567452), (43195,-0.724393), (43196,-0.744309), (43197,-0.924938), (43198,-0.922557), (43199,-1.069285), (43200,-1.176058), (43201,-0.935858), (43202,-0.638064), (43203,-0.811723), (43204,-0.872986), (43205,-0.938419), (43206,-0.764180), (43207,-0.908579), (43208,-0.879723), (43209,-0.620012), (43210,-0.342656), (43211,-0.499134), (43212,-0.558994), (43213,-0.744269), (43214,-0.734461), (43215,-0.917876), (43216,-0.981919), (43217,-0.729647), (43218,-0.466217), (43219,-0.601793), (43220,-0.639361), (43221,-0.698295), (43222,-0.537061), (43223,-0.694929), (43224,-1.013985), (43225,-0.769139), (43226,-0.497349), (43227,-0.636645), (43228,-0.729948), (43229,-0.898041), (43230,-0.864076), (43231,-1.004292), (43232,-1.047903), (43233,-0.851360), (43234,-0.561462), (43235,-0.716543), (43236,-0.815426), (43237,-0.871109), (43238,-0.698260), (43239,-0.853811), (43240,-0.878837), (43241,-0.543880), (43242,-0.684096), (43243,-0.413703), (43244,-0.590155), (43245,-0.683928), (43246,-0.857124), (43247,-0.821769), (43248,-0.962918), (43249,-0.640966), (43250,-0.783975), (43251,-0.489431), (43252,-0.612928), (43253,-0.609620), (43254,-0.771207), (43255,-0.643411), (43256,-0.707923), (43257,-0.856035), (43258,-0.174570), (43259,-0.324541), (43260,-0.387657), (43261,-0.567359), (43262,-0.598422), (43263,-0.785093), (43264,-0.719081), (43265,-0.910862), (43266,-0.234499), (43267,-0.404446), (43268,-0.439691), (43269,-0.615210), (43270,-0.395912), (43271,-0.492472), (43272,-0.695862), (43273,-0.735290), (43274,-0.531784), (43275,-0.268823), (43276,-0.444349), (43277,-0.498173), (43278,-0.655577), (43279,-0.625331), (43280,-0.789705), (43281,-0.858394), (43282,-0.613078), (43283,-0.318534), (43284,-0.466652), (43285,-0.514903), (43286,-0.558971), (43287,-0.424212), (43288,-0.797143), (43289,-0.513281), (43290,-0.323244), (43291,-0.353379), (43292,-0.503821), (43293,-0.485184), (43294,-0.660710), (43295,-0.699668), (43296,-0.871474), (43297,-0.567174), (43298,-0.328828), (43299,-0.366397), (43300,-0.548422), (43301,-0.362104), (43302,-0.440085), (43303,-0.508768), (43304,-0.856621), (43305,-0.624318), (43306,-0.338132), (43307,-0.489964), (43308,-0.540074), (43309,-0.696088), (43310,-0.696030), (43311,-0.844612), (43312,-0.897509), (43313,-0.671705), (43314,-0.374838), (43315,-0.554076), (43316,-0.611613), (43317,-0.679375), (43318,-0.540897), (43319,-0.695521), (43320,-0.785575), (43321,-0.527723), (43322,-0.289841), (43323,-0.345988), (43324,-0.515477), (43325,-0.474543), (43326,-0.666787), (43327,-0.744298), (43328,-0.897990), (43329,-0.608555), (43330,-0.366495), (43331,-0.409637), (43332,-0.560541), (43333,-0.378863), (43334,-0.453595), (43335,-0.505096), (43336,-0.675042), (43337,-0.833379), (43338,-0.172809), (43339,-0.280984), (43340,-0.320869), (43341,-0.491285), (43342,-0.512592), (43343,-0.694617), (43344,-0.756806), (43345,-0.897028), (43346,-0.227629), (43347,-0.395258), (43348,-0.460698), (43349,-0.631571), (43350,-0.332380), (43351,-0.478175), (43352,-0.749385), (43353,-0.501284), (43354,-0.232750), (43355,-0.276824), (43356,-0.437478), (43357,-0.410946), (43358,-0.626878), (43359,-0.672343), (43360,-0.826497), (43361,-0.529166), (43362,-0.287107), (43363,-0.379484), (43364,-0.511810), (43365,-0.349644), (43366,-0.418332), (43367,-0.433603), (43368,-0.735470), (43369,-0.489228), (43370,-0.238810), (43371,-0.438950), (43372,-0.476518), (43373,-0.660403), (43374,-0.630151), (43375,-0.786166), (43376,-0.858568), (43377,-0.625338), (43378,-0.314531), (43379,-0.458004), (43380,-0.506254), (43381,-0.556828), (43382,-0.439257), (43383,-0.574827), (43384,-0.906425), (43385,-0.602125), (43386,-0.354956), (43387,-0.475204), (43388,-0.539246), (43389,-0.701760), (43390,-0.742115), (43391,-0.899519), (43392,-1.188844), (43393,-0.539889), (43394,-0.690331), (43395,-0.743228), (43396,-0.887626), (43397,-0.650677), (43398,-0.818770), (43399,-0.845186), (43400,-0.899943), (43401,-0.683894), (43402,-0.380984), (43403,-0.589954), (43404,-0.619156), (43405,-0.775634), (43406,-0.791374), (43407,-0.945992), (43408,-1.010498), (43409,-0.757293), (43410,-0.458102), (43411,-0.621086), (43412,-0.680946), (43413,-0.779828), (43414,-0.610693), (43415,-0.788072), (43416,-1.019332), (43417,-0.761018), (43418,-0.504563), (43419,-0.659644), (43420,-0.734839), (43421,-0.899676), (43422,-0.888472), (43423,-1.050523), (43424,-1.098773), (43425,-0.916639), (43426,-0.583535), (43427,-0.731653), (43428,-0.758075), (43429,-0.826758), (43430,-0.699432), (43431,-0.824789), (43432,-0.925525), (43433,-0.674179), (43434,-0.427474), (43435,-0.576989), (43436,-0.609441), (43437,-0.750127), (43438,-0.783519), (43439,-0.917235), (43440,-0.980351), (43441,-0.741078), (43442,-0.460003), (43443,-0.642491), (43444,-0.675414), (43445,-0.751535), (43446,-0.580540), (43447,-0.732377), (43448,-1.057000), (43449,-0.800075), (43450,-0.524579), (43451,-0.699171), (43452,-0.755781), (43453,-0.910863), (43454,-0.919633), (43455,-1.101659), (43456,-1.116003), (43457,-0.877193), (43458,-0.628634), (43459,-0.740516), (43460,-0.804565), (43461,-0.906228), (43462,-0.739885), (43463,-0.915868), (43464,-0.900024), (43465,-0.703481), (43466,-0.392681), (43467,-0.541726), (43468,-0.586258), (43469,-0.771069), (43470,-0.757542), (43471,-0.918666), (43472,-0.948338), (43473,-0.703029), (43474,-0.405699), (43475,-0.573322), (43476,-0.650370), (43477,-0.731601), (43478,-0.550393), (43479,-0.759819), (43480,-1.056577), (43481,-0.784324), (43482,-0.514864), (43483,-0.688060), (43484,-0.740494), (43485,-0.898831), (43486,-0.851391), (43487,-1.015301), (43488,-1.110001), (43489,-0.826139), (43490,-0.557605), (43491,-0.708046), (43492,-0.754438), (43493,-0.832882), (43494,-0.681861), (43495,-0.875965), (43496,-0.934899), (43497,-0.694699), (43498,-0.395045), (43499,-0.553376), (43500,-0.616955), (43501,-0.817096), (43502,-0.792886), (43503,-0.944718), (43504,-0.985536), (43505,-0.756952), (43506,-0.456365), (43507,-0.594264), (43508,-0.668526), (43509,-0.711204), (43510,-0.572725), (43511,-0.719453), (43512,-0.702670), (43513,-0.873086), (43514,-0.216699), (43515,-0.345769), (43516,-0.410745), (43517,-0.579764), (43518,-0.594571), (43519,-0.762195), (43520,-0.778392), (43521,-0.932553), (43522,-0.298920), (43523,-0.413131), (43524,-0.506441), (43525,-0.685210), (43526,-0.433865), (43527,-0.606134), (43528,-0.779800), (43529,-0.943241), (43530,-0.232044), (43531,-0.410820), (43532,-0.499483), (43533,-0.679649), (43534,-0.661939), (43535,-0.791942), (43536,-0.835547), (43537,-0.976696), (43538,-0.269213), (43539,-0.423374), (43540,-0.486947), (43541,-0.615090), (43542,-0.397189), (43543,-0.538801), (43544,-0.829516), (43545,-0.541014), (43546,-0.318460), (43547,-0.377393), (43548,-0.513903), (43549,-0.526850), (43550,-0.675432), (43551,-0.756663), (43552,-0.893165), (43553,-0.637174), (43554,-0.398828), (43555,-0.441969), (43556,-0.603093), (43557,-0.455792), (43558,-0.560247), (43559,-0.605712), (43560,-1.048316), (43561,-0.321792), (43562,-0.463404), (43563,-0.554854), (43564,-0.686247), (43565,-0.701518), (43566,-0.880293), (43567,-0.909966), (43568,-1.066443), (43569,-0.415628), (43570,-0.534016), (43571,-0.572981), (43572,-0.751287), (43573,-0.503654), (43574,-0.641554), (43575,-0.674939), (43576,-0.797046), (43577,-0.469522), (43578,-0.292027), (43579,-0.351423), (43580,-0.496292), (43581,-0.501807), (43582,-0.675009), (43583,-0.722790), (43584,-0.869982), (43585,-0.620027), (43586,-0.384004), (43587,-0.458735), (43588,-0.590128), (43589,-0.427498), (43590,-0.505010), (43591,-0.553261), (43592,-0.791027), (43593,-0.515525), (43594,-0.281362), (43595,-0.342618), (43596,-0.496772), (43597,-0.474423), (43598,-0.652728), (43599,-0.680078), (43600,-0.856067), (43601,-0.568485), (43602,-0.343614), (43603,-0.363531), (43604,-0.534874), (43605,-0.399651), (43606,-0.469730), (43607,-0.544925), (43608,-0.776649), (43609,-0.468166), (43610,-0.205206), (43611,-0.283650), (43612,-0.433622), (43613,-0.438210), (43614,-0.625814), (43615,-0.679638), (43616,-0.846798), (43617,-0.575941), (43618,-0.326913), (43619,-0.392815), (43620,-0.535824), (43621,-0.382017), (43622,-0.473930), (43623,-0.554235), (43624,-0.870961), (43625,-0.189952), (43626,-0.333424), (43627,-0.372852), (43628,-0.504709), (43629,-0.504188), (43630,-0.677390), (43631,-0.751652), (43632,-0.941573), (43633,-0.280076), (43634,-0.409616), (43635,-0.465299), (43636,-0.606911), (43637,-0.389003), (43638,-0.521330), (43639,-0.558898), (43640,-1.008472), (43641,-0.316781), (43642,-0.493696), (43643,-0.545197), (43644,-0.673347), (43645,-0.732280), (43646,-0.894794), (43647,-0.963019), (43648,-1.014983), (43649,-0.747377), (43650,-0.486276), (43651,-0.639040), (43652,-0.720265), (43653,-0.789423), (43654,-0.602173), (43655,-0.773515), (43656,-0.940675), (43657,-0.691647), (43658,-0.425436), (43659,-0.565659), (43660,-0.630165), (43661,-0.827055), (43662,-0.807492), (43663,-0.962573), (43664,-0.982953), (43665,-0.775734), (43666,-0.508127), (43667,-0.631161), (43668,-0.680808), (43669,-0.771789), (43670,-0.584075), (43671,-0.761460), (43672,-0.903536), (43673,-0.570438), (43674,-0.733885), (43675,-0.451876), (43676,-0.599068), (43677,-0.666824), (43678,-0.823301), (43679,-0.861333), (43680,-1.037322), (43681,-0.669384), (43682,-0.814716), (43683,-0.564761), (43684,-0.743067), (43685,-0.692846), (43686,-0.817740), (43687,-0.703882), (43688,-0.699178), (43689,-0.727924), (43690,-0.885792), (43691,-0.575919), (43692,-0.756084), (43693,-0.799689), (43694,-0.959886), (43695,-0.966797), (43696,-0.730311), (43697,-0.774379), (43698,-0.934112), (43699,-0.690193), (43700,-0.737048), (43701,-0.813633), (43702,-1.011456), (43703,-0.838137), (43704,-1.014590), (43705,-0.642476), (43706,-0.775265), (43707,-0.528097), (43708,-0.685964), (43709,-0.737471), (43710,-0.885583), (43711,-0.885995), (43712,-1.053618), (43713,-0.718661), (43714,-0.859810), (43715,-0.580130), (43716,-0.679940), (43717,-0.643188), (43718,-0.817318), (43719,-0.657004), (43720,-0.858541), (43721,-0.539839), (43722,-0.679598), (43723,-0.391090), (43724,-0.580547), (43725,-0.668278), (43726,-0.804781), (43727,-0.800546), (43728,-0.927293), (43729,-0.590483), (43730,-0.741387), (43731,-0.450093), (43732,-0.620502), (43733,-0.589324), (43734,-0.752307), (43735,-0.604073), (43736,-0.938921), (43737,-0.617432), (43738,-0.743716), (43739,-0.484475), (43740,-0.627014), (43741,-0.703599), (43742,-0.833602), (43743,-0.812642), (43744,-0.936140), (43745,-0.611871), (43746,-0.766489), (43747,-0.480767), (43748,-0.655823), (43749,-0.627901), (43750,-0.778805), (43751,-0.660765), (43752,-0.840467), (43753,-0.488321), (43754,-0.602996), (43755,-0.340499), (43756,-0.465392), (43757,-0.557306), (43758,-0.695668), (43759,-0.684464), (43760,-0.867880), (43761,-0.492046), (43762,-0.630409), (43763,-0.385563), (43764,-0.518822), (43765,-0.442121), (43766,-0.614854), (43767,-0.478705), (43768,-0.765701), (43769,-0.453041), (43770,-0.570966), (43771,-0.316365), (43772,-0.444045), (43773,-0.491832), (43774,-0.678503), (43775,-0.710029), (43776,-0.837246), (43777,-0.518081), (43778,-0.636005), (43779,-0.361435), (43780,-0.495152), (43781,-0.471406), (43782,-0.642749), (43783,-0.521922), (43784,-0.820996), (43785,-0.496258), (43786,-0.648559), (43787,-0.355868), (43788,-0.471933), (43789,-0.582431), (43790,-0.747268), (43791,-0.722595), (43792,-0.906010), (43793,-0.567803), (43794,-0.737286), (43795,-0.460857), (43796,-0.594110), (43797,-0.545279), (43798,-0.712903), (43799,-0.547023), (43800,-0.801972), (43801,-0.595679), (43802,-0.332719), (43803,-0.465508), (43804,-0.515155), (43805,-0.718082), (43806,-0.736602), (43807,-0.878221), (43808,-0.919039), (43809,-0.652359), (43810,-0.367570), (43811,-0.512432), (43812,-0.553251), (43813,-0.647951), (43814,-0.518764), (43815,-0.666883), (43816,-0.751363), (43817,-0.552967), (43818,-0.242167), (43819,-0.380530), (43820,-0.434353), (43821,-0.607549), (43822,-0.594023), (43823,-0.748647), (43824,-0.806647), (43825,-0.558551), (43826,-0.311852), (43827,-0.453928), (43828,-0.513325), (43829,-0.601062), (43830,-0.449114), (43831,-0.601409), (43832,-0.834529), (43833,-0.576215), (43834,-0.293280), (43835,-0.460903), (43836,-0.492898), (43837,-0.681429), (43838,-0.678122), (43839,-0.826233), (43840,-0.877740), (43841,-0.661229), (43842,-0.367611), (43843,-0.553349), (43844,-0.604387), (43845,-0.657284), (43846,-0.501623), (43847,-0.703617), (43848,-0.837803), (43849,-0.600853), (43850,-0.311418), (43851,-0.478115), (43852,-0.534261), (43853,-0.698172), (43854,-0.686961), (43855,-0.820684), (43856,-0.902379), (43857,-0.689580), (43858,-0.429869), (43859,-0.534788), (43860,-0.600691), (43861,-0.659161), (43862,-0.549949), (43863,-0.705963), (43864,-0.842466), (43865,-0.620845), (43866,-0.298430), (43867,-0.485101), (43868,-0.514774), (43869,-0.678677), (43870,-0.684199), (43871,-0.834640), (43872,-0.855483), (43873,-0.615284), (43874,-0.352787), (43875,-0.526916), (43876,-0.593745), (43877,-0.650355), (43878,-0.469147), (43879,-0.612156), (43880,-0.526632), (43881,-0.680323), (43882,-0.377876), (43883,-0.521348), (43884,-0.590037), (43885,-0.765100), (43886,-0.742744), (43887,-0.893185), (43888,-0.572160), (43889,-0.715632), (43890,-0.412258), (43891,-0.540872), (43892,-0.539417), (43893,-0.686145), (43894,-0.547203), (43895,-0.710650), (43896,-0.773297), (43897,-0.542390), (43898,-0.220901), (43899,-0.389921), (43900,-0.477651), (43901,-0.635989), (43902,-0.615492), (43903,-0.803554), (43904,-1.095202), (43905,-0.750952), (43906,-0.916259), (43907,-0.616605), (43908,-0.733133), (43909,-0.684303), (43910,-0.903028), (43911,-0.757580), (43912,-1.019034), (43913,-0.701265), (43914,-0.833585), (43915,-0.512103), (43916,-0.710384), (43917,-0.800437), (43918,-0.956452), (43919,-0.975905), (43920,-1.109158), (43921,-0.766305), (43922,-0.893985), (43923,-0.628238), (43924,-0.785179), (43925,-0.783261), (43926,-0.892363), (43927,-0.745061), (43928,-0.860199), (43929,-0.898694), (43930,-0.707730), (43931,-0.418759), (43932,-0.569664), (43933,-0.625347), (43934,-0.790647), (43935,-0.769224), (43936,-0.903874), (43937,-0.921931), (43938,-0.726321), (43939,-0.446635), (43940,-0.581284), (43941,-0.647187), (43942,-0.718662), (43943,-0.556032), (43944,-0.786830), (43945,-0.590756), (43946,-0.681737), (43947,-0.824745), (43948,-0.502794), (43949,-0.668563), (43950,-0.732606), (43951,-0.896516), (43952,-0.875557), (43953,-0.656722), (43954,-0.696614), (43955,-0.843799), (43956,-0.618928), (43957,-0.695513), (43958,-0.744690), (43959,-0.863085), (43960,-1.058115), (43961,-0.719902), (43962,-0.870806), (43963,-0.586944), (43964,-0.716484), (43965,-0.818153), (43966,-0.951870), (43967,-0.959708), (43968,-1.125941), (43969,-0.777978), (43970,-0.936779), (43971,-0.673355), (43972,-0.834942), (43973,-0.799117), (43974,-0.955595), (43975,-0.816189), (43976,-0.940150), (43977,-0.660471), (43978,-0.763067), (43979,-0.905612), (43980,-0.576227), (43981,-0.772648), (43982,-0.872927), (43983,-1.041941), (43984,-1.012622), (43985,-0.792397), (43986,-0.835538), (43987,-0.974828), (43988,-0.714190), (43989,-0.801457), (43990,-0.827880), (43991,-0.948128), (43992,-0.945283), (43993,-0.967059), (43994,-0.754724), (43995,-0.466680), (43996,-0.622694), (43997,-0.630068), (43998,-0.856689), (43999,-0.837583), (44000,-0.969909), (44001,-1.013051), (44002,-0.756126), (44003,-0.496885), (44004,-0.678447), (44005,-0.716479), (44006,-0.779588), (44007,-0.582588), (44008,-0.696800), (44009,-0.880678), (44010,-0.515064), (44011,-0.675724), (44012,-0.403941), (44013,-0.523725), (44014,-0.596127), (44015,-0.735416), (44016,-0.781807), (44017,-0.938291), (44018,-0.597755), (44019,-0.734264), (44020,-0.474089), (44021,-0.630104), (44022,-0.637015), (44023,-0.780017), (44024,-0.778569), (44025,-0.821247), (44026,-0.539238), (44027,-0.258163), (44028,-0.425329), (44029,-0.473574), (44030,-0.624015), (44031,-0.614207), (44032,-0.768362), (44033,-0.771554), (44034,-0.562938), (44035,-0.297654), (44036,-0.397464), (44037,-0.465689), (44038,-0.581760), (44039,-0.405655), (44040,-0.608119), (44041,-0.752987), (44042,-0.456120), (44043,-0.584726), (44044,-0.294358), (44045,-0.426685), (44046,-0.510232), (44047,-0.661607), (44048,-0.648543), (44049,-0.810594), (44050,-0.490032), (44051,-0.608426), (44052,-0.376586), (44053,-0.526558), (44054,-0.521396), (44055,-0.654649), (44056,-0.819950), (44057,-0.880742), (44058,-0.613599), (44059,-0.322768), (44060,-0.508049), (44061,-0.564196), (44062,-0.724850), (44063,-0.710396), (44064,-0.865014), (44065,-0.954604), (44066,-0.738093), (44067,-0.446798), (44068,-0.584697), (44069,-0.643630), (44070,-0.730434), (44071,-0.574774), (44072,-0.791169), (44073,-0.829664), (44074,-0.580642), (44075,-0.277269), (44076,-0.420278), (44077,-0.469455), (44078,-0.663096), (44079,-0.637490), (44080,-0.755878), (44081,-0.860333), (44082,-0.600623), (44083,-0.317693), (44084,-0.453733), (44085,-0.508947), (44086,-0.546978), (44087,-0.424761), (44088,-0.740098), (44089,-0.791135), (44090,-0.571374), (44091,-0.244776), (44092,-0.419368), (44093,-0.454613), (44094,-0.674265), (44095,-0.649123), (44096,-0.820465), (44097,-0.858034), (44098,-0.589031), (44099,-0.330253), (44100,-0.503919), (44101,-0.528945), (44102,-0.586945), (44103,-0.470301), (44104,-0.728506), (44105,-0.778616), (44106,-0.570001), (44107,-0.273133), (44108,-0.427751), (44109,-0.448131), (44110,-0.623650), (44111,-0.614306), (44112,-0.773570), (44113,-0.806956), (44114,-0.599273), (44115,-0.297760), (44116,-0.446341), (44117,-0.518280), (44118,-0.586042), (44119,-0.431308), (44120,-0.771259), (44121,-0.854813), (44122,-0.597425), (44123,-0.314027), (44124,-0.489082), (44125,-0.545693), (44126,-0.741656), (44127,-0.705368), (44128,-0.866955), (44129,-0.916596), (44130,-0.700085), (44131,-0.388821), (44132,-0.530897), (44133,-0.593550), (44134,-0.670598), (44135,-0.493566), (44136,-0.765703), (44137,-0.445148), (44138,-0.597442), (44139,-0.361426), (44140,-0.523940), (44141,-0.637218), (44142,-0.761185), (44143,-0.752768), (44144,-0.932006), (44145,-0.593329), (44146,-0.749344), (44147,-0.420892), (44148,-0.593162), (44149,-0.544332), (44150,-0.698486), (44151,-0.579519), (44152,-0.951523), (44153,-0.593341), (44154,-0.708943), (44155,-0.444122), (44156,-0.614075), (44157,-0.673471), (44158,-0.852710), (44159,-0.848469), (44160,-1.234412), (44161,-0.918960), (44162,-1.066151), (44163,-0.771137), (44164,-0.948516), (44165,-0.927563), (44166,-1.075675), (44167,-0.942776), (44168,-1.172177), (44169,-0.814458), (44170,-0.957467), (44171,-0.691256), (44172,-0.824509), (44173,-0.897381), (44174,-1.099838), (44175,-1.089104), (44176,-1.227930), (44177,-0.866492), (44178,-1.041554), (44179,-0.718206), (44180,-0.896055), (44181,-0.854187), (44182,-1.009275), (44183,-0.865687), (44184,-1.036103), (44185,-1.088530), (44186,-0.822320), (44187,-0.520343), (44188,-0.680533), (44189,-0.741326), (44190,-0.921961), (44191,-0.940482), (44192,-1.083027), (44193,-1.143357), (44194,-0.889219), (44195,-0.606747), (44196,-0.741396), (44197,-0.819371), (44198,-0.875518), (44199,-0.698956), (44200,-1.013365), (44201,-0.776879), (44202,-0.838135), (44203,-0.979747), (44204,-0.687526), (44205,-0.886733), (44206,-0.970287), (44207,-1.084962), (44208,-1.075148), (44209,-0.810798), (44210,-0.856725), (44211,-1.024812), (44212,-0.753029), (44213,-0.819858), (44214,-0.888547), (44215,-1.069175), (44216,-1.213117), (44217,-0.872117), (44218,-1.017912), (44219,-0.749842), (44220,-0.888668), (44221,-0.973619), (44222,-1.083647), (44223,-1.101241), (44224,-1.251212), (44225,-0.913005), (44226,-1.061587), (44227,-0.777261), (44228,-0.927696), (44229,-0.896055), (44230,-1.053928), (44231,-0.922882), (44232,-0.975779), (44233,-0.732794), (44234,-0.795903), (44235,-0.959350), (44236,-0.658763), (44237,-0.861226), (44238,-0.908087), (44239,-1.055272), (44240,-1.051964), (44241,-0.804796), (44242,-0.876741), (44243,-1.048077), (44244,-0.765148), (44245,-0.845910), (44246,-0.924354), (44247,-1.031596), (44248,-1.059872), (44249,-1.069570), (44250,-0.866064), (44251,-0.552471), (44252,-0.696876), (44253,-0.748377), (44254,-0.936438), (44255,-0.910369), (44256,-1.071030), (44257,-1.120207), (44258,-0.899056), (44259,-0.624016), (44260,-0.799072), (44261,-0.838037), (44262,-0.897897), (44263,-0.745023), (44264,-0.801170), (44265,-0.925600), (44266,-0.593429), (44267,-0.795892), (44268,-0.497165), (44269,-0.637844), (44270,-0.725581), (44271,-0.836073), (44272,-0.800712), (44273,-1.003175), (44274,-0.629665), (44275,-0.797758), (44276,-0.517145), (44277,-0.664800), (44278,-0.629902), (44279,-0.769661), (44280,-0.783072), (44281,-0.846188), (44282,-0.598556), (44283,-0.330022), (44284,-0.485573), (44285,-0.488765), (44286,-0.702374), (44287,-0.717645), (44288,-0.880628), (44289,-0.915410), (44290,-0.664058), (44291,-0.403421), (44292,-0.584983), (44293,-0.619765), (44294,-0.689380), (44295,-0.529537), (44296,-0.762194), (44297,-0.923318), (44298,-0.596720), (44299,-0.733686), (44300,-0.473981), (44301,-0.634172), (44302,-0.716793), (44303,-0.849583), (44304,-0.812368), (44305,-0.957230), (44306,-0.628779), (44307,-0.777824), (44308,-0.533441), (44309,-0.653689), (44310,-0.625766), (44311,-0.802682), (44312,-0.938721), (44313,-1.021343), (44314,-0.783003), (44315,-0.470337), (44316,-0.661191), (44317,-0.685284), (44318,-0.840372), (44319,-0.844960), (44320,-0.974494), (44321,-1.040859), (44322,-0.782082), (44323,-0.519584), (44324,-0.667703), (44325,-0.710381), (44326,-0.779996), (44327,-0.617366), (44328,-0.814257), (44329,-0.888518), (44330,-0.616265), (44331,-0.364920), (44332,-0.515362), (44333,-0.565929), (44334,-0.754924), (44335,-0.736287), (44336,-0.861644), (44337,-0.906182), (44338,-0.686884), (44339,-0.416021), (44340,-0.594333), (44341,-0.670455), (44342,-0.756325), (44343,-0.594629), (44344,-0.841218), (44345,-0.855562), (44346,-0.611643), (44347,-0.363547), (44348,-0.484722), (44349,-0.523680), (44350,-0.730790), (44351,-0.724695), (44352,-0.894178), (44353,-0.940106), (44354,-0.695724), (44355,-0.416971), (44356,-0.602253), (44357,-0.639815), (44358,-0.728478), (44359,-0.552843), (44360,-0.820797), (44361,-0.912710), (44362,-0.662292), (44363,-0.398405), (44364,-0.540480), (44365,-0.597097), (44366,-0.761934), (44367,-0.770698), (44368,-0.941578), (44369,-0.966141), (44370,-0.694351), (44371,-0.402593), (44372,-0.555821), (44373,-0.618937), (44374,-0.695985), (44375,-0.540324), (44376,-0.910932), (44377,-0.935959), (44378,-0.686930), (44379,-0.425829), (44380,-0.594849), (44381,-0.644490), (44382,-0.789358), (44383,-0.749820), (44384,-0.925803), (44385,-1.013077), (44386,-0.766835), (44387,-0.485296), (44388,-0.662211), (44389,-0.685841), (44390,-0.801912), (44391,-0.638813), (44392,-0.984806), (44393,-0.603400), (44394,-0.733403), (44395,-0.482984), (44396,-0.643638), (44397,-0.742058), (44398,-0.898999), (44399,-0.898014), (44400,-1.036376), (44401,-0.681908), (44402,-0.840708), (44403,-0.549414), (44404,-0.665948), (44405,-0.709089), (44406,-0.853951), (44407,-0.676926), (44408,-1.021060), (44409,-0.680060), (44410,-0.861158), (44411,-0.559181), (44412,-0.701257), (44413,-0.770409), (44414,-0.933856), (44415,-0.931475), (44416,-1.069374), (44417,-1.124131), (44418,-0.883461), (44419,-0.602849), (44420,-0.768619), (44421,-0.803401), (44422,-0.886022), (44423,-0.718746), (44424,-0.969518), (44425,-1.022878), (44426,-0.778960), (44427,-0.490921), (44428,-0.664117), (44429,-0.707722), (44430,-0.850267), (44431,-0.830234), (44432,-1.009010), (44433,-1.077699), (44434,-0.843072), (44435,-0.541095), (44436,-0.677598), (44437,-0.731421), (44438,-0.820085), (44439,-0.655596), (44440,-1.010881), (44441,-1.056809), (44442,-0.868168), (44443,-0.584769), (44444,-0.760752), (44445,-0.772773), (44446,-0.926927), (44447,-0.918047), (44448,-1.124223), (44449,-1.179443), (44450,-0.939244), (44451,-0.631694), (44452,-0.777019), (44453,-0.841995), (44454,-0.906038), (44455,-0.721573), (44456,-0.808377), (44457,-0.945813), (44458,-0.626184), (44459,-0.789168), (44460,-0.547109), (44461,-0.704976), (44462,-0.830797), (44463,-0.940362), (44464,-0.915689), (44465,-1.016425), (44466,-0.676822), (44467,-0.831446), (44468,-0.594033), (44469,-0.716603), (44470,-0.717935), (44471,-0.858621), (44472,-1.003953), (44473,-1.015510), (44474,-0.767878), (44475,-0.489589), (44476,-0.690656), (44477,-0.749589), (44478,-0.922792), (44479,-0.927380), (44480,-1.081534), (44481,-1.129322), (44482,-0.881220), (44483,-0.608973), (44484,-0.731544), (44485,-0.819274), (44486,-0.882390), (44487,-0.730443), (44488,-0.814924), (44489,-0.966292), (44490,-0.627152), (44491,-0.757155), (44492,-0.479799), (44493,-0.686902), (44494,-0.753731), (44495,-0.873052), (44496,-0.833977), (44497,-0.986742), (44498,-0.652711), (44499,-0.824981), (44500,-0.566666), (44501,-0.718498), (44502,-0.688252), (44503,-0.818719), (44504,-1.010030), (44505,-1.076396), (44506,-0.846879), (44507,-0.555121), (44508,-0.729250), (44509,-0.824413), (44510,-0.996219), (44511,-1.009167), (44512,-1.163327), (44513,-1.224114), (44514,-0.977878), (44515,-0.675438), (44516,-0.834238), (44517,-0.879696), (44518,-0.926557), (44519,-0.787615), (44520,-0.848872), (44521,-1.006276), (44522,-0.656460), (44523,-0.808754), (44524,-0.537434), (44525,-0.641427), (44526,-0.737053), (44527,-0.872166), (44528,-0.837268), (44529,-0.988173), (44530,-0.639283), (44531,-0.794828), (44532,-0.573213), (44533,-0.678132), (44534,-0.643234), (44535,-0.795998), (44536,-0.805696), (44537,-0.894823), (44538,-0.651831), (44539,-0.367969), (44540,-0.559749), (44541,-0.618683), (44542,-0.777483), (44543,-0.755134), (44544,-0.845187), (44545,-0.904584), (44546,-0.680176), (44547,-0.369377), (44548,-0.546756), (44549,-0.622877), (44550,-0.710608), (44551,-0.557734), (44552,-0.769020), (44553,-0.925034), (44554,-0.566852), (44555,-0.738658), (44556,-0.431572), (44557,-0.579683), (44558,-0.670207), (44559,-0.822501), (44560,-0.802012), (44561,-0.943161), (44562,-0.651866), (44563,-0.783723), (44564,-0.479886), (44565,-0.653552), (44566,-0.637702), (44567,-0.746803), (44568,-0.734667), (44569,-0.789423), (44570,-0.911061), (44571,-0.245387), (44572,-0.381427), (44573,-0.440823), (44574,-0.591728), (44575,-0.585170), (44576,-0.789950), (44577,-0.835878), (44578,-1.033701), (44579,-0.335041), (44580,-0.483159), (44581,-0.522581), (44582,-0.664200), (44583,-0.429573), (44584,-0.843844), (44585,-0.916246), (44586,-0.650499), (44587,-0.388471), (44588,-0.583502), (44589,-0.621997), (44590,-0.786370), (44591,-0.787245), (44592,-0.928394), (44593,-0.969212), (44594,-0.710898), (44595,-0.467442), (44596,-0.623920), (44597,-0.698182), (44598,-0.749682), (44599,-0.577766), (44600,-0.843867), (44601,-0.878179), (44602,-0.650985), (44603,-0.344362), (44604,-0.505949), (44605,-0.581607), (44606,-0.739938), (44607,-0.740350), (44608,-0.920052), (44609,-0.993387), (44610,-0.749468), (44611,-0.476752), (44612,-0.635553), (44613,-0.700992), (44614,-0.745993), (44615,-0.594045), (44616,-0.846671), (44617,-0.875410), (44618,-0.646363), (44619,-0.371323), (44620,-0.518509), (44621,-0.522633), (44622,-0.691190), (44623,-0.698564), (44624,-0.901954), (44625,-0.975289), (44626,-0.763424), (44627,-0.492567), (44628,-0.657868), (44629,-0.705192), (44630,-0.747870), (44631,-0.572698), (44632,-0.697122), (44633,-0.755592), (44634,-0.879559), (44635,-0.218061), (44636,-0.384758), (44637,-0.444618), (44638,-0.584377), (44639,-0.597787), (44640,-0.765417), (44641,-0.824350), (44642,-0.954817), (44643,-0.306325), (44644,-0.425639), (44645,-0.502224), (44646,-0.608540), (44647,-0.367877), (44648,-0.753350), (44649,-0.832721), (44650,-0.581840), (44651,-0.307727), (44652,-0.473960), (44653,-0.537539), (44654,-0.722814), (44655,-0.687459), (44656,-0.850900), (44657,-0.902407), (44658,-0.682639), (44659,-0.417825), (44660,-0.559901), (44661,-0.598866), (44662,-0.605307), (44663,-0.470548), (44664,-0.809572), (44665,-0.871292), (44666,-0.630629), (44667,-0.364882), (44668,-0.535292), (44669,-0.570537), (44670,-0.757208), (44671,-0.696769), (44672,-1.119862), (44673,-0.753784), (44674,-0.939066), (44675,-0.658917), (44676,-0.824217), (44677,-0.768424), (44678,-0.929084), (44679,-0.782710), (44680,-0.912713), (44681,-0.713853), (44682,-0.774640), (44683,-0.935300), (44684,-0.658407), (44685,-0.826957), (44686,-0.877531), (44687,-1.016357), (44688,-1.019092), (44689,-0.786318), (44690,-0.807632), (44691,-0.960859), (44692,-0.689070), (44693,-0.794922), (44694,-0.814369), (44695,-0.998254), (44696,-0.823082), (44697,-0.954481), (44698,-0.620451), (44699,-0.792720), (44700,-0.534869), (44701,-0.664409), (44702,-0.736348), (44703,-0.906294), (44704,-0.872329), (44705,-1.060397), (44706,-0.724043), (44707,-0.859619), (44708,-0.588299), (44709,-0.753599), (44710,-0.736359), (44711,-0.847314), (44712,-0.994969), (44713,-0.780781), (44714,-0.823453), (44715,-0.965535), (44716,-0.690032), (44717,-0.828394), (44718,-0.896150), (44719,-1.036836), (44720,-1.050716), (44721,-0.807730), (44722,-0.849475), (44723,-1.030110), (44724,-0.751821), (44725,-0.820973), (44726,-0.869224), (44727,-1.005264), (44728,-1.050728), (44729,-0.771975), (44730,-0.852737), (44731,-0.967411), (44732,-0.691445), (44733,-0.864642), (44734,-0.918935), (44735,-1.063797), (44736,-1.038198), (44737,-0.794742), (44738,-0.892228), (44739,-1.028738), (44740,-0.714218), (44741,-0.803339), (44742,-0.846017), (44743,-1.019683), (44744,-0.910008), (44745,-0.648901), (44746,-0.711553), (44747,-0.865245), (44748,-0.580913), (44749,-0.747609), (44750,-0.788434), (44751,-0.948625), (44752,-0.910477), (44753,-0.711154), (44754,-0.758941), (44755,-0.957685), (44756,-0.650598), (44757,-0.713714), (44758,-0.771257), (44759,-0.904974), (44760,-0.798549), (44761,-0.970355), (44762,-0.603344), (44763,-0.749139), (44764,-0.493148), (44765,-0.650089), (44766,-0.712741), (44767,-0.834842), (44768,-0.891459), (44769,-1.056295), (44770,-0.703223), (44771,-0.856914), (44772,-0.576765), (44773,-0.730920), (44774,-0.680699), (44775,-0.865048), (44776,-0.716813), (44777,-0.831951), (44778,-0.501640), (44779,-0.675769), (44780,-0.393297), (44781,-0.520514), (44782,-0.598959), (44783,-0.735462), (44784,-0.753055), (44785,-0.916039), (44786,-0.534632), (44787,-0.693896), (44788,-0.416997), (44789,-0.611564), (44790,-0.568777), (44791,-0.713176), (44792,-0.690826), (44793,-0.779020), (44794,-0.438026), (44795,-0.633984), (44796,-0.339439), (44797,-0.484771), (44798,-0.522339), (44799,-0.692749), (44800,-0.628127), (44801,-0.783678), (44802,-0.440361), (44803,-0.610771), (44804,-0.394259), (44805,-0.545627), (44806,-0.484255), (44807,-0.635630), (44808,-0.624889), (44809,-0.756746), (44810,-0.439440), (44811,-0.600100), (44812,-0.366401), (44813,-0.528914), (44814,-0.612932), (44815,-0.789847), (44816,-0.755882), (44817,-0.890068), (44818,-0.574616), (44819,-0.720411), (44820,-0.447232), (44821,-0.587454), (44822,-0.540020), (44823,-0.695565), (44824,-0.888272), (44825,-0.942102), (44826,-0.674032), (44827,-0.378555), (44828,-0.568476), (44829,-0.618586), (44830,-0.790392), (44831,-0.791724), (44832,-0.960744), (44833,-1.011318), (44834,-0.792483), (44835,-0.474714), (44836,-0.629802), (44837,-0.688735), (44838,-0.732340), (44839,-0.584575), (44840,-0.723401), (44841,-0.741921), (44842,-0.513801), (44843,-0.279637), (44844,-0.442151), (44845,-0.524779), (44846,-0.676147), (44847,-0.672839), (44848,-0.821420), (44849,-0.869671), (44850,-0.640617), (44851,-0.358609), (44852,-0.527165), (44853,-0.569843), (44854,-0.608338), (44855,-0.465683), (44856,-0.744789), (44857,-0.791180), (44858,-0.593247), (44859,-0.301952), (44860,-0.458430), (44861,-0.487639), (44862,-0.654799), (44863,-0.613865), (44864,-0.828407), (44865,-0.860866), (44866,-0.606264), (44867,-0.315433), (44868,-0.510000), (44869,-0.557324), (44870,-0.593033), (44871,-0.459664), (44872,-0.686279), (44873,-0.718274), (44874,-0.478075), (44875,-0.223010), (44876,-0.363232), (44877,-0.401264), (44878,-0.616263), (44879,-0.590664), (44880,-0.763397), (44881,-0.839055), (44882,-0.572838), (44883,-0.319633), (44884,-0.481220), (44885,-0.539227), (44886,-0.659011), (44887,-0.454578), (44888,-0.823790), (44889,-0.912917), (44890,-0.669467), (44891,-0.395355), (44892,-0.535114), (44893,-0.593120), (44894,-0.764926), (44895,-0.748143), (44896,-0.885579), (44897,-0.938476), (44898,-0.686661), (44899,-0.387934), (44900,-0.579715), (44901,-0.647007), (44902,-0.712910), (44903,-0.586510), (44904,-0.849824), (44905,-0.615661), (44906,-0.659266), (44907,-0.746533), (44908,-0.477073), (44909,-0.656775), (44910,-0.733823), (44911,-0.862430), (44912,-0.835897), (44913,-0.596161), (44914,-0.653705), (44915,-0.775805), (44916,-0.526320), (44917,-0.612191), (44918,-0.687849), (44919,-0.877307), (44920,-0.933917), (44921,-0.612428), (44922,-0.778662), (44923,-0.497586), (44924,-0.632235), (44925,-0.683736), (44926,-0.821635), (44927,-0.814145), (44928,-0.542825), (44929,-0.302625), (44930,-0.369918), (44931,-0.535688), (44932,-0.250892), (44933,-0.319581), (44934,-0.384557), (44935,-0.529419), (44936,-0.486162), (44937,-0.251535), (44938,-0.280281), (44939,-0.419570), (44940,-0.167762), (44941,-0.370219), (44942,-0.416153), (44943,-0.548936), (44944,-0.567926), (44945,-0.372779), (44946,-0.395483), (44947,-0.549174), (44948,-0.240697), (44949,-0.273619), (44950,-0.381325), (44951,-0.526187), (44952,-0.483862), (44953,-0.238090), (44954,-0.304456), (44955,-0.420057), (44956,-0.155700), (44957,-0.327506), (44958,-0.390159), (44959,-0.560105), (44960,-0.548902), (44961,-0.304983), (44962,-0.350447), (44963,-0.520400), (44964,-0.248610), (44965,-0.321945), (44966,-0.376232), (44967,-0.524814), (44968,-0.235379), (44969,-0.323573), (44970,-0.480983), (44971,-0.511583), (44972,-0.686175), (44973,-0.373516), (44974,-0.552285), (44975,-0.580567), (44976,-0.339898), (44977,-0.326834), (44978,-0.483782), (44979,-0.541782), (44980,-0.614654), (44981,-0.341474), (44982,-0.472404), (44983,-0.533197), (44984,-0.506664), (44985,-0.302232), (44986,-0.363488), (44987,-0.504173), (44988,-0.211019), (44989,-0.419519), (44990,-0.451977), (44991,-0.600096), (44992,-0.621402), (44993,-0.359838), (44994,-0.434100), (44995,-0.585931), (44996,-0.274662), (44997,-0.367972), (44998,-0.419009), (44999,-0.603357), (45000,-0.400315), (45001,-0.082076), (45002,-0.221835), (45003,-0.309102), (45004,-0.464190), (45005,-0.202156), (45006,-0.355383), (45007,-0.413390), (45008,-0.567081), (45009,-0.139219), (45010,-0.313348), (45011,-0.394579), (45012,-0.552917), (45013,-0.174297), (45014,-0.336810), (45015,-0.378098), (45016,-0.527143), (45017,-0.259073), (45018,-0.303141), (45019,-0.467051), (45020,-0.181329), (45021,-0.376823), (45022,-0.432507), (45023,-0.595490), (45024,-0.569421), (45025,-0.303674), (45026,-0.346352), (45027,-0.504220), (45028,-0.213858), (45029,-0.302515), (45030,-0.334974), (45031,-0.449649), (45032,-0.324645), (45033,-0.007803), (45034,-0.159171), (45035,-0.189307), (45036,-0.359253), (45037,-0.126950), (45038,-0.256483), (45039,-0.325636), (45040,-0.476540), (45041,-0.054727), (45042,-0.238606), (45043,-0.301722), (45044,-0.456803), (45045,-0.081903), (45046,-0.268574), (45047,-0.309392), (45048,-0.405019), (45049,-0.172252), (45050,-0.224216), (45051,-0.355615), (45052,-0.087545), (45053,-0.251919), (45054,-0.328967), (45055,-0.495200), (45056,-0.441724), (45057,-0.214067), (45058,-0.266031), (45059,-0.400217), (45060,-0.137256), (45061,-0.224060), (45062,-0.287170), (45063,-0.426465), (45064,-0.436163), (45065,-0.125357), (45066,-0.299949), (45067,-0.337518), (45068,-0.481916), (45069,-0.220815), (45070,-0.352209), (45071,-0.416721), (45072,-0.548114), (45073,-0.137911), (45074,-0.300888), (45075,-0.354248), (45076,-0.484715), (45077,-0.099595), (45078,-0.233775), (45079,-0.326152), (45080,-0.379512), (45081,-0.128630), (45082,-0.181990), (45083,-0.346364), (45084,-0.081543), (45085,-0.289580), (45086,-0.351769), (45087,-0.524502), (45088,-0.510975), (45089,-0.268452), (45090,-0.266541), (45091,-0.397001), (45092,-0.092701), (45093,-0.221778), (45094,-0.263986), (45095,-0.425573), (45096,-0.333086), (45097,-0.062230), (45098,-0.113730), (45099,-0.255806), (45100,0.000649), (45101,-0.177194), (45102,-0.237523), (45103,-0.402823), (45104,-0.390230), (45105,-0.163499), (45106,-0.200598), (45107,-0.342680), (45108,-0.043952), (45109,-0.140042), (45110,-0.189690), (45111,-0.367068), (45112,-0.430648), (45113,-0.221569), (45114,-0.238699), (45115,-0.378452), (45116,-0.108992), (45117,-0.262683), (45118,-0.339268), (45119,-0.494818), (45120,-0.471073), (45121,-0.217398), (45122,-0.293519), (45123,-0.495983), (45124,-0.198182), (45125,-0.291955), (45126,-0.330914), (45127,-0.449308), (45128,-0.413483), (45129,-0.193722), (45130,-0.206669), (45131,-0.364073), (45132,-0.052341), (45133,-0.254804), (45134,-0.301665), (45135,-0.453959), (45136,-0.429287), (45137,-0.186301), (45138,-0.223863), (45139,-0.379877), (45140,-0.119703), (45141,-0.205117), (45142,-0.247325), (45143,-0.418668), (45144,-0.366588), (45145,-0.133821), (45146,-0.205296), (45147,-0.332977), (45148,-0.059334), (45149,-0.245072), (45150,-0.282177), (45151,-0.408924), (45152,-0.392147), (45153,-0.155198), (45154,-0.190443), (45155,-0.358530), (45156,-0.070021), (45157,-0.178660), (45158,-0.210655), (45159,-0.352731), (45160,-0.014987), (45161,-0.199335), (45162,-0.274987), (45163,-0.418929), (45164,-0.141103), (45165,-0.317086), (45166,-0.366733), (45167,-0.499986), (45168,-0.154810), (45169,-0.297355), (45170,-0.311229), (45171,-0.502547), (45172,-0.154584), (45173,-0.301306), (45174,-0.359312), (45175,-0.489779), (45176,-0.367092), (45177,-0.124106), (45178,-0.169571), (45179,-0.336267), (45180,-0.078879), (45181,-0.241863), (45182,-0.269676), (45183,-0.426616), (45184,-0.515743), (45185,-0.167317), (45186,-0.325185), (45187,-0.209004), (45188,-0.373847), (45189,-0.358461), (45190,-0.486141), (45191,-0.209705), (45192,-0.469306), (45193,-0.148281), (45194,-0.288967), (45195,-0.289835), (45196,-0.447709), (45197,-0.496887), (45198,-0.627817), (45199,-0.383904), (45200,-0.553387), (45201,-0.222613), (45202,-0.371194), (45203,-0.214137), (45204,-0.345067), (45205,-0.305060), (45206,-0.460610), (45207,-0.179071), (45208,-0.420088), (45209,-0.175706), (45210,-0.235102), (45211,-0.417127), (45212,-0.363194), (45213,-0.566120), (45214,-0.622267), (45215,-0.784318), (45216,-0.494413), (45217,-0.236562), (45218,-0.281563), (45219,-0.481703), (45220,-0.320470), (45221,-0.388226), (45222,-0.410002), (45223,-0.597137), (45224,-0.370406), (45225,-0.094903), (45226,-0.125503), (45227,-0.273621), (45228,-0.321408), (45229,-0.495537), (45230,-0.535892), (45231,-0.679364), (45232,-0.434049), (45233,-0.200819), (45234,-0.242564), (45235,-0.387895), (45236,-0.228985), (45237,-0.290241), (45238,-0.369613), (45239,-0.511688), (45240,-0.367174), (45241,-0.113042), (45242,-0.166402), (45243,-0.352604), (45244,-0.347436), (45245,-0.490445), (45246,-0.535446), (45247,-0.694710), (45248,-0.432676), (45249,-0.199909), (45250,-0.279281), (45251,-0.382810), (45252,-0.238758), (45253,-0.318593), (45254,-0.377063), (45255,-0.531680), (45256,-0.298450), (45257,-0.061964), (45258,-0.090240), (45259,-0.239755), (45260,-0.212759), (45261,-0.413362), (45262,-0.495983), (45263,-0.617627), (45264,-0.325863), (45265,-0.080554), (45266,-0.147383), (45267,-0.327092), (45268,-0.158419), (45269,-0.249406), (45270,-0.288364), (45271,-0.461567), (45272,-0.409950), (45273,-0.184610), (45274,-0.223111), (45275,-0.398167), (45276,-0.369775), (45277,-0.579671), (45278,-0.599124), (45279,-0.753742), (45280,-0.504714), (45281,-0.238967), (45282,-0.307655), (45283,-0.474815), (45284,-0.340056), (45285,-0.405959), (45286,-0.468611), (45287,-0.609760), (45288,-0.375134), (45289,-0.153976), (45290,-0.207336), (45291,-0.354991), (45292,-0.369329), (45293,-0.529063), (45294,-0.535974), (45295,-0.716603), (45296,-0.448069), (45297,-0.217156), (45298,-0.262157), (45299,-0.429317), (45300,-0.254145), (45301,-0.295896), (45302,-0.341360), (45303,-0.496441), (45304,-0.253455), (45305,-0.017433), (45306,-0.091231), (45307,-0.207302), (45308,-0.202598), (45309,-0.394842), (45310,-0.458885), (45311,-0.626508), (45312,-0.377486), (45313,-0.103380), (45314,-0.163239), (45315,-0.325753), (45316,-0.176599), (45317,-0.221593), (45318,-0.272630), (45319,-0.414712), (45320,-0.330579), (45321,-0.113141), (45322,-0.149782), (45323,-0.303473), (45324,-0.298769), (45325,-0.476612), (45326,-0.480736), (45327,-0.619099), (45328,-0.338950), (45329,-0.088532), (45330,-0.154434), (45331,-0.283041), (45332,-0.165007), (45333,-0.239268), (45334,-0.305171), (45335,-0.502518), (45336,-0.275794), (45337,-0.324972), (45338,-0.044359), (45339,-0.048484), (45340,-0.210071), (45341,-0.287119), (45342,-0.461712), (45343,-0.145803), (45344,-0.299024), (45345,-0.364000), (45346,-0.122867), (45347,0.037439), (45348,-0.142726), (45349,-0.192373), (45350,-0.263849), (45351,0.048348), (45352,-0.390074), (45353,-0.080201), (45354,-0.220423), (45355,-0.232444), (45356,-0.370807), (45357,-0.448782), (45358,-0.564853), (45359,-0.299569), (45360,-0.462083), (45361,-0.159179), (45362,-0.278493), (45363,-0.109827), (45364,-0.278384), (45365,-0.254638), (45366,-0.406469), (45367,-0.123070), (45368,-0.388238), (45369,-0.070006), (45370,-0.186070), (45371,-0.214346), (45372,-0.358282), (45373,-0.444622), (45374,-0.611782), (45375,-0.323280), (45376,-0.475112), (45377,-0.129935), (45378,-0.280840), (45379,-0.166982), (45380,-0.318350), (45381,-0.274630), (45382,-0.397664), (45383,-0.115192), (45384,-0.366890), (45385,-0.081175), (45386,-0.246475), (45387,-0.224589), (45388,-0.377817), (45389,-0.391228), (45390,-0.557924), (45391,-0.288458), (45392,-0.476062), (45393,-0.116484), (45394,-0.292473), (45395,-0.160963), (45396,-0.322087), (45397,-0.281616), (45398,-0.432521), (45399,-0.103600), (45400,-0.231743), (45401,-0.248874), (45402,-0.021216), (45403,-0.004440), (45404,-0.175313), (45405,-0.212881), (45406,-0.397229), (45407,-0.124513), (45408,-0.288423), (45409,-0.393342), (45410,-0.139674), (45411,0.013200), (45412,-0.132589), (45413,-0.172480), (45414,-0.239779), (45415,0.054309), (45416,-0.289825), (45417,0.032590), (45418,-0.131783), (45419,-0.111294), (45420,-0.259405), (45421,-0.345283), (45422,-0.508729), (45423,-0.232763), (45424,-0.373449), (45425,-0.061716), (45426,-0.212151), (45427,-0.035589), (45428,-0.210182), (45429,-0.185509), (45430,-0.339200), (45431,-0.030717), (45432,-0.344194), (45433,-0.009236), (45434,-0.148526), (45435,-0.134999), (45436,-0.306805), (45437,-0.413583), (45438,-0.569598), (45439,-0.313606), (45440,-0.457542), (45441,-0.225238), (45442,-0.263270), (45443,-0.376548), (45444,-0.249685), (45445,-0.322087), (45446,-0.404245), (45447,-0.575588), (45448,-0.387873), (45449,-0.107731), (45450,-0.160158), (45451,-0.327324), (45452,-0.304969), (45453,-0.499536), (45454,-0.581694), (45455,-0.720989), (45456,-0.451523), (45457,-0.209464), (45458,-0.247495), (45459,-0.426734), (45460,-0.272463), (45461,-0.334183), (45462,-0.389403), (45463,-0.535662), (45464,-0.736265), (45465,-0.066872), (45466,-0.222423), (45467,-0.274387), (45468,-0.410432), (45469,-0.433136), (45470,-0.587290), (45471,-0.638791), (45472,-0.780403), (45473,-0.125875), (45474,-0.284212), (45475,-0.342682), (45476,-0.504732), (45477,-0.278929), (45478,-0.450271), (45479,-0.477621), (45480,-0.651287), (45481,-0.011617), (45482,-0.162985), (45483,-0.182902), (45484,-0.358891), (45485,-0.343968), (45486,-0.489300), (45487,-0.549629), (45488,-0.718185), (45489,-0.031604), (45490,-0.183435), (45491,-0.245155), (45492,-0.400242), (45493,-0.128922), (45494,-0.289576), (45495,-0.349443), (45496,-0.700076), (45497,0.006474), (45498,-0.163472), (45499,-0.222869), (45500,-0.351945), (45501,-0.377898), (45502,-0.531589), (45503,-0.584023), (45504,-0.727032), (45505,-0.055315), (45506,-0.234084), (45507,-0.291164), (45508,-0.438349), (45509,-0.200936), (45510,-0.344408), (45511,-0.419597), (45512,-0.624853), (45513,0.100282), (45514,-0.046440), (45515,-0.092831), (45516,-0.263711), (45517,-0.293383), (45518,-0.439641), (45519,-0.479063), (45520,-0.640187), (45521,0.025487), (45522,-0.132844), (45523,-0.198283), (45524,-0.389131), (45525,-0.124317), (45526,-0.294263), (45527,-0.336941), (45528,-0.737280), (45529,-0.050235), (45530,-0.204389), (45531,-0.301412), (45532,-0.454640), (45533,-0.439253), (45534,-0.597591), (45535,-0.642585), (45536,-0.810215), (45537,-0.097159), (45538,-0.244808), (45539,-0.336258), (45540,-0.459292), (45541,-0.220019), (45542,-0.411336), (45543,-0.490708), (45544,-0.643009), (45545,0.068194), (45546,-0.119874), (45547,-0.183917), (45548,-0.317633), (45549,-0.339873), (45550,-0.470803), (45551,-0.559466), (45552,-0.716871), (45553,-0.060483), (45554,-0.198382), (45555,-0.272644), (45556,-0.431444), (45557,-0.162448), (45558,-0.357009), (45559,-0.432203), (45560,-0.481381), (45561,-0.200305), (45562,0.032925), (45563,-0.008357), (45564,-0.146719), (45565,-0.106718), (45566,-0.326363), (45567,-0.377400), (45568,-0.569181), (45569,-0.321086), (45570,-0.035364), (45571,-0.093371), (45572,-0.232660), (45573,-0.063061), (45574,-0.128037), (45575,-0.171641), (45576,-0.459570), (45577,-0.206365), (45578,0.013860), (45579,-0.037178), (45580,-0.180650), (45581,-0.167123), (45582,-0.364940), (45583,-0.435019), (45584,-0.577101), (45585,-0.283483), (45586,-0.071618), (45587,-0.113363), (45588,-0.288882), (45589,-0.140191), (45590,-0.201910), (45591,-0.257130), (45592,-0.173460), (45593,-0.316005), (45594,0.032884), (45595,-0.089680), (45596,-0.092878), (45597,-0.254002), (45598,-0.320368), (45599,-0.446188), (45600,-0.222707), (45601,-0.377795), (45602,-0.020540), (45603,-0.155652), (45604,-0.022283), (45605,-0.235429), (45606,-0.207970), (45607,-0.331931), (45608,-0.356957), (45609,-0.083314), (45610,-0.164545), (45611,-0.316840), (45612,-0.315392), (45613,-0.475582), (45614,-0.528016), (45615,-0.648727), (45616,-0.346750), (45617,-0.176687), (45618,-0.244449), (45619,-0.422292), (45620,-0.271277), (45621,-0.310699), (45622,-0.332476), (45623,-0.467582), (45624,-0.142380), (45625,-0.314186), (45626,0.009619), (45627,-0.131994), (45628,-0.131935), (45629,-0.305601), (45630,-0.404014), (45631,-0.519152), (45632,-0.233900), (45633,-0.380622), (45634,-0.031726), (45635,-0.138042), (45636,-0.035330), (45637,-0.193667), (45638,-0.158312), (45639,-0.314320), (45640,-0.134045), (45641,-0.296558), (45642,0.050478), (45643,-0.100427), (45644,-0.093869), (45645,-0.294009), (45646,-0.344583), (45647,-0.491305), (45648,-0.212553), (45649,-0.392255), (45650,-0.049865), (45651,-0.197520), (45652,-0.053932), (45653,-0.196007), (45654,-0.178304), (45655,-0.331532), (45656,-0.127092), (45657,-0.285893), (45658,0.015157), (45659,-0.122279), (45660,-0.114788), (45661,-0.255010), (45662,-0.328809), (45663,-0.512694), (45664,-0.224649), (45665,-0.367657), (45666,0.000744), (45667,-0.146442), (45668,0.005969), (45669,-0.178842), (45670,-0.118403), (45671,-0.266985), (45672,-0.196326), (45673,0.042020), (45674,-0.028529), (45675,-0.165965), (45676,-0.137109), (45677,-0.327030), (45678,-0.341368), (45679,-0.513644), (45680,-0.207484), (45681,0.015997), (45682,-0.055942), (45683,-0.216139), (45684,-0.111567), (45685,-0.192798), (45686,-0.207605), (45687,-0.346431), (45688,-0.238146), (45689,-0.002593), (45690,-0.088470), (45691,-0.227296), (45692,-0.186362), (45693,-0.374423), (45694,-0.421284), (45695,-0.542458), (45696,-0.536364), (45697,-0.306847), (45698,-0.364390), (45699,-0.500893), (45700,-0.383316), (45701,-0.433890), (45702,-0.492823), (45703,-0.628869), (45704,-0.426753), (45705,-0.189340), (45706,-0.257102), (45707,-0.447023), (45708,-0.425600), (45709,-0.605766), (45710,-0.637761), (45711,-0.790056), (45712,-0.488542), (45713,-0.251593), (45714,-0.314245), (45715,-0.467467), (45716,-0.318775), (45717,-0.388391), (45718,-0.430142), (45719,-0.612167), (45720,-0.654376), (45721,-0.372373), (45722,-0.140533), (45723,-0.201789), (45724,-0.313678), (45725,-0.291322), (45726,-0.482639), (45727,-0.501623), (45728,-0.675752), (45729,-0.415578), (45730,-0.188384), (45731,-0.236635), (45732,-0.413550), (45733,-0.245811), (45734,-0.274557), (45735,-0.332557), (45736,-0.644180), (45737,-0.015193), (45738,-0.134977), (45739,-0.224104), (45740,-0.348998), (45741,-0.380524), (45742,-0.514710), (45743,-0.592685), (45744,-0.727798), (45745,-0.033783), (45746,-0.159604), (45747,-0.248731), (45748,-0.388490), (45749,-0.198453), (45750,-0.360503), (45751,-0.436161), (45752,-0.797946), (45753,-0.120194), (45754,-0.272025), (45755,-0.356969), (45756,-0.519020), (45757,-0.551479), (45758,-0.681482), (45759,-0.731123), (45760,-0.902935), (45761,-0.216817), (45762,-0.355643), (45763,-0.434551), (45764,-0.571987), (45765,-0.393565), (45766,-0.522635), (45767,-0.578318), (45768,-0.752448), (45769,-0.034746), (45770,-0.208411), (45771,-0.256192), (45772,-0.392702), (45773,-0.414941), (45774,-0.571419), (45775,-0.628492), (45776,-0.828169), (45777,-0.152270), (45778,-0.290633), (45779,-0.350962), (45780,-0.484678), (45781,-0.251912), (45782,-0.416285), (45783,-0.476615), (45784,-0.671182), (45785,-0.382674), (45786,-0.126213), (45787,-0.187006), (45788,-0.336984), (45789,-0.325774), (45790,-0.480861), (45791,-0.520283), (45792,-0.648896), (45793,-0.392435), (45794,-0.168491), (45795,-0.193517), (45796,-0.348141), (45797,-0.239393), (45798,-0.312258), (45799,-0.350290), (45800,-0.543931), (45801,-0.250776), (45802,-0.029619), (45803,-0.084839), (45804,-0.202300), (45805,-0.213851), (45806,-0.402845), (45807,-0.444127), (45808,-0.578776), (45809,-0.285622), (45810,-0.078403), (45811,-0.140122), (45812,-0.253864), (45813,-0.091704), (45814,-0.165966), (45815,-0.233258), (45816,-0.402278), (45817,-0.165791), (45818,0.091596), (45819,0.033590), (45820,-0.140539), (45821,-0.133982), (45822,-0.283027), (45823,-0.321522), (45824,-0.528631), (45825,-0.227581), (45826,0.026087), (45827,-0.065826), (45828,-0.180964), (45829,-0.036449), (45830,-0.109315), (45831,-0.191942), (45832,-0.519814), (45833,-0.239202), (45834,-0.005972), (45835,-0.033784), (45836,-0.169824), (45837,-0.170229), (45838,-0.325317), (45839,-0.368458), (45840,-0.512857), (45841,-0.265688), (45842,-0.034317), (45843,-0.118798), (45844,-0.261337), (45845,-0.122402), (45846,-0.159037), (45847,-0.263029), (45848,-0.193761), (45849,-0.323764), (45850,0.046033), (45851,-0.129023), (45852,-0.140580), (45853,-0.318423), (45854,-0.348558), (45855,-0.511542), (45856,-0.247185), (45857,-0.404595), (45858,-0.035261), (45859,-0.197318), (45860,-0.081601), (45861,-0.232505), (45862,-0.181352), (45863,-0.361054), (45864,-0.227691), (45865,-0.360944), (45866,-0.019945), (45867,-0.167136), (45868,-0.139671), (45869,-0.298471), (45870,-0.377379), (45871,-0.551045), (45872,-0.273683), (45873,-0.448275), (45874,-0.133756), (45875,-0.301386), (45876,-0.128537), (45877,-0.285478), (45878,-0.281237), (45879,-0.412173), (45880,-0.225849), (45881,-0.345170), (45882,-0.005566), (45883,-0.197347), (45884,-0.215404), (45885,-0.374668), (45886,-0.402017), (45887,-0.544099), (45888,-0.295998), (45889,-0.457585), (45890,-0.098940), (45891,-0.249381), (45892,-0.067240), (45893,-0.283641), (45894,-0.209264), (45895,-0.371777), (45896,-0.203575), (45897,-0.352620), (45898,-0.020449), (45899,-0.184829), (45900,-0.198703), (45901,-0.339852), (45902,-0.418296), (45903,-0.562695), (45904,-0.286266), (45905,-0.400007), (45906,-0.045081), (45907,-0.200626), (45908,-0.047752), (45909,-0.233496), (45910,-0.195812), (45911,-0.365758), (45912,-0.156216), (45913,-0.327559), (45914,-0.007003), (45915,-0.134214), (45916,-0.133692), (45917,-0.296676), (45918,-0.363968), (45919,-0.575724), (45920,-0.259808), (45921,-0.406067), (45922,-0.034416), (45923,-0.174638), (45924,-0.020368), (45925,-0.190778), (45926,-0.174934), (45927,-0.301681), (45928,-0.244492), (45929,-0.030303), (45930,-0.093419), (45931,-0.267079), (45932,-0.258661), (45933,-0.438363), (45934,-0.493120), (45935,-0.637519), (45936,-0.368985), (45937,-0.129713), (45938,-0.176573), (45939,-0.316326), (45940,-0.168561), (45941,-0.253975), (45942,-0.291537), (45943,-0.457771), (45944,-0.459572), (45945,-0.212867), (45946,-0.274123), (45947,-0.434784), (45948,-0.395709), (45949,-0.580984), (45950,-0.648283), (45951,-0.816370), (45952,-0.524148), (45953,-0.639286), (45954,-0.296433), (45955,-0.456624), (45956,-0.311645), (45957,-0.459764), (45958,-0.448096), (45959,-0.574844), (45960,-0.721565), (45961,-0.446996), (45962,-0.183108), (45963,-0.215098), (45964,-0.395263), (45965,-0.421222), (45966,-0.592095), (45967,-0.630127), (45968,-0.775459), (45969,-0.457690), (45970,-0.218880), (45971,-0.243907), (45972,-0.391098), (45973,-0.269338), (45974,-0.335704), (45975,-0.381638), (45976,-0.652842), (45977,-0.369907), (45978,-0.093941), (45979,-0.210938), (45980,-0.362306), (45981,-0.334847), (45982,-0.533128), (45983,-0.550721), (45984,-0.706272), (45985,-0.445165), (45986,-0.210538), (45987,-0.262972), (45988,-0.430595), (45989,-0.258679), (45990,-0.359879), (45991,-0.419745), (45992,-0.832626), (45993,-0.153940), (45994,-0.318314), (45995,-0.359595), (45996,-0.451045), (45997,-0.488150), (45998,-0.679461), (45999,-0.752796), (46000,-0.878617), (46001,-0.215729), (46002,-0.393572), (46003,-0.427890), (46004,-0.556961), (46005,-0.319084), (46006,-0.468593), (46007,-0.524739), (46008,-0.743928), (46009,-0.467028), (46010,-0.201281), (46011,-0.214692), (46012,-0.401364), (46013,-0.382727), (46014,-0.546637), (46015,-0.569340), (46016,-0.765767), (46017,-0.510239), (46018,-0.229627), (46019,-0.289487), (46020,-0.460367), (46021,-0.317711), (46022,-0.370602), (46023,-0.422572), (46024,-0.632468), (46025,-0.385300), (46026,-0.141381), (46027,-0.188241), (46028,-0.344256), (46029,-0.317254), (46030,-0.517857), (46031,-0.589802), (46032,-0.690538), (46033,-0.406676), (46034,-0.170190), (46035,-0.218904), (46036,-0.380491), (46037,-0.260597), (46038,-0.322780), (46039,-0.381250), (46040,-0.658496), (46041,-0.391359), (46042,-0.146977), (46043,-0.230995), (46044,-0.395831), (46045,-0.394383), (46046,-0.542965), (46047,-0.619086), (46048,-0.775564), (46049,-0.505171), (46050,-0.247320), (46051,-0.287674), (46052,-0.446938), (46053,-0.273626), (46054,-0.327450), (46055,-0.406821), (46056,-0.576304), (46057,-0.297552), (46058,-0.052706), (46059,-0.096311), (46060,-0.246752), (46061,-0.319154), (46062,-0.504429), (46063,-0.496475), (46064,-0.636697), (46065,-0.349116), (46066,-0.127031), (46067,-0.137662), (46068,-0.314114), (46069,-0.170526), (46070,-0.252221), (46071,-0.316727), (46072,-0.641355), (46073,-0.338908), (46074,-0.063875), (46075,-0.117699), (46076,-0.271390), (46077,-0.254607), (46078,-0.422700), (46079,-0.489066), (46080,-0.623246), (46081,-0.349603), (46082,-0.101971), (46083,-0.185525), (46084,-0.313205), (46085,-0.186342), (46086,-0.259670), (46087,-0.328359), (46088,-0.646945), (46089,-0.328713), (46090,-0.101519), (46091,-0.145124), (46092,-0.292309), (46093,-0.305726), (46094,-0.474276), (46095,-0.552721), (46096,-0.688760), (46097,-0.398398), (46098,-0.136828), (46099,-0.210163), (46100,-0.357348), (46101,-0.195182), (46102,-0.297784), (46103,-0.332559), (46104,-0.294881), (46105,-0.441140), (46106,-0.122438), (46107,-0.294244), (46108,-0.263998), (46109,-0.386099), (46110,-0.478013), (46111,-0.647032), (46112,-0.367816), (46113,-0.478308), (46114,-0.128022), (46115,-0.336058), (46116,-0.179002), (46117,-0.342448), (46118,-0.284332), (46119,-0.449632), (46120,-0.201537), (46121,-0.309706), (46122,0.004814), (46123,-0.155383), (46124,-0.148356), (46125,-0.291365), (46126,-0.403253), (46127,-0.562980), (46128,-0.288874), (46129,-0.436523), (46130,-0.072768), (46131,-0.205094), (46132,-0.053610), (46133,-0.230989), (46134,-0.194238), (46135,-0.345606), (46136,-0.280520), (46137,-0.431425), (46138,-0.106223), (46139,-0.243189), (46140,-0.221766), (46141,-0.376854), (46142,-0.486419), (46143,-0.615489), (46144,-0.371107), (46145,-0.543846), (46146,-0.215388), (46147,-0.339819), (46148,-0.204127), (46149,-0.344812), (46150,-0.296445), (46151,-0.438527), (46152,-0.254063), (46153,-0.398468), (46154,-0.061188), (46155,-0.216269), (46156,-0.209248), (46157,-0.357829), (46158,-0.425585), (46159,-0.585782), (46160,-0.336291), (46161,-0.475580), (46162,-0.137373), (46163,-0.258084), (46164,-0.118215), (46165,-0.270979), (46166,-0.235618), (46167,-0.370267), (46168,-0.167225), (46169,-0.314416), (46170,0.021011), (46171,-0.144759), (46172,-0.148420), (46173,-0.287710), (46174,-0.347576), (46175,-0.523095), (46176,-0.281963), (46177,-0.469567), (46178,-0.111385), (46179,-0.272503), (46180,-0.127988), (46181,-0.283539), (46182,-0.283481), (46183,-0.428812), (46184,-0.351648), (46185,-0.090084), (46186,-0.148554), (46187,-0.321287), (46188,-0.273389), (46189,-0.471207), (46190,-0.534323), (46191,-0.694513), (46192,-0.427370), (46193,-0.171842), (46194,-0.225665), (46195,-0.395155), (46196,-0.212550), (46197,-0.289598), (46198,-0.347605), (46199,-0.549605), (46200,-0.290357), (46201,-0.409208), (46202,-0.090049), (46203,-0.227016), (46204,-0.217672), (46205,-0.387155), (46206,-0.482318), (46207,-0.612321), (46208,-0.758579), (46209,-0.512337), (46210,-0.243804), (46211,-0.288342), (46212,-0.430881), (46213,-0.295195), (46214,-0.380602), (46215,-0.453004), (46216,-0.692167), (46217,-0.430597), (46218,-0.180178), (46219,-0.231679), (46220,-0.380261), (46221,-0.368130), (46222,-0.542723), (46223,-0.609552), (46224,-0.756274), (46225,-0.463589), (46226,-0.235925), (46227,-0.299505), (46228,-0.453665), (46229,-0.306828), (46230,-0.356468), (46231,-0.390324), (46232,-0.733061), (46233,-0.445016), (46234,-0.225718), (46235,-0.271182), (46236,-0.460640), (46237,-0.437358), (46238,-0.610560), (46239,-0.677389), (46240,-0.838976), (46241,-0.560224), (46242,-0.315841), (46243,-0.357586), (46244,-0.512674), (46245,-0.348648), (46246,-0.407117), (46247,-0.431217), (46248,-0.757699), (46249,-0.107817), (46250,-0.263362), (46251,-0.329727), (46252,-0.481095), (46253,-0.514487), (46254,-0.651917), (46255,-0.715033), (46256,-0.876620), (46257,-0.216049), (46258,-0.389252), (46259,-0.469550), (46260,-0.594443), (46261,-0.375146), (46262,-0.506075), (46263,-0.570118), (46264,-0.780014), (46265,-0.496615), (46266,-0.210430), (46267,-0.267510), (46268,-0.410512), (46269,-0.405351), (46270,-0.579480), (46271,-0.661638), (46272,-0.825548), (46273,-0.530071), (46274,-0.296371), (46275,-0.326043), (46276,-0.501099), (46277,-0.327324), (46278,-0.430383), (46279,-0.453556), (46280,-0.685743), (46281,-0.374474), (46282,-0.134274), (46283,-0.150478), (46284,-0.341789), (46285,-0.346377), (46286,-0.547914), (46287,-0.602664), (46288,-0.758678), (46289,-0.461811), (46290,-0.240653), (46291,-0.304696), (46292,-0.456997), (46293,-0.269746), (46294,-0.332862), (46295,-0.373217), (46296,-0.744288), (46297,-0.460426), (46298,-0.222086), (46299,-0.303781), (46300,-0.439357), (46301,-0.412355), (46302,-0.567442), (46303,-0.640777), (46304,-0.824656), (46305,-0.567738), (46306,-0.300131), (46307,-0.377643), (46308,-0.535517), (46309,-0.381246), (46310,-0.480592), (46311,-0.514441), (46312,-0.556656), (46313,-0.698268), (46314,-0.020979), (46315,-0.189535), (46316,-0.239639), (46317,-0.409129), (46318,-0.393279), (46319,-0.534428), (46320,-0.603116), (46321,-0.775386), (46322,-0.090201), (46323,-0.229490), (46324,-0.290746), (46325,-0.482527), (46326,-0.232109), (46327,-0.373721), (46328,-0.580367), (46329,-0.262592), (46330,-0.034471), (46331,-0.100837), (46332,-0.274033), (46333,-0.250750), (46334,-0.415594), (46335,-0.454552), (46336,-0.617072), (46337,-0.355038), (46338,-0.081395), (46339,-0.151474), (46340,-0.296343), (46341,-0.125347), (46342,-0.213547), (46343,-0.253902), (46344,-0.450323), (46345,-0.631885), (46346,0.058873), (46347,-0.094818), (46348,-0.145855), (46349,-0.335313), (46350,-0.369625), (46351,-0.503811), (46352,-0.565067), (46353,-0.698320), (46354,-0.022885), (46355,-0.156138), (46356,-0.249447), (46357,-0.393383), (46358,-0.148537), (46359,-0.273431), (46360,-0.097332), (46361,-0.249164), (46362,-0.279763), (46363,-0.035381), (46364,-0.001879), (46365,-0.189947), (46366,-0.264672), (46367,-0.431368), (46368,-0.129391), (46369,-0.311416), (46370,-0.374996), (46371,-0.147802), (46372,0.010651), (46373,-0.154655), (46374,-0.208015), (46375,-0.266022), (46376,-0.578565), (46377,-0.314215), (46378,-0.067973), (46379,-0.134338), (46380,-0.293139), (46381,-0.250351), (46382,-0.433303), (46383,-0.468549), (46384,-0.682621), (46385,-0.375071), (46386,-0.139981), (46387,-0.161758), (46388,-0.354002), (46389,-0.186726), (46390,-0.264237), (46391,-0.311561), (46392,-0.246939), (46393,-0.395984), (46394,-0.070319), (46395,-0.232833), (46396,-0.218843), (46397,-0.358132), (46398,-0.409169), (46399,-0.567970), (46400,-0.304083), (46401,-0.450341), (46402,-0.120493), (46403,-0.260246), (46404,-0.106445), (46405,-0.261990), (46406,-0.253572), (46407,-0.403550), (46408,-0.543772), (46409,-0.258514), (46410,-0.045716), (46411,-0.072138), (46412,-0.190526), (46413,-0.219272), (46414,-0.402687), (46415,-0.440255), (46416,-0.593483), (46417,-0.311011), (46418,-0.078244), (46419,-0.129281), (46420,-0.307124), (46421,-0.169115), (46422,-0.267065), (46423,-0.288841), (46424,-0.091371), (46425,-0.272470), (46426,-0.297959), (46427,-0.096776), (46428,-0.047019), (46429,-0.193741), (46430,-0.268936), (46431,-0.470466), (46432,-0.194500), (46433,-0.363057), (46434,-0.375077), (46435,-0.122799), (46436,0.021716), (46437,-0.142194), (46438,-0.190445), (46439,-0.266097), (46440,-0.665509), (46441,-0.029096), (46442,-0.202755), (46443,-0.244970), (46444,-0.397271), (46445,-0.381884), (46446,-0.523497), (46447,-0.595435), (46448,-0.709647), (46449,-0.035607), (46450,-0.196267), (46451,-0.252414), (46452,-0.403319), (46453,-0.222574), (46454,-0.367899), (46455,-0.456563), (46456,-0.627443), (46457,-0.359836), (46458,-0.130782), (46459,-0.163241), (46460,-0.306250), (46461,-0.272748), (46462,-0.450127), (46463,-0.509524), (46464,-0.723602), (46465,-0.444380), (46466,-0.204181), (46467,-0.259401), (46468,-0.374539), (46469,-0.231414), (46470,-0.315901), (46471,-0.375761), (46472,-0.657654), (46473,-0.358463), (46474,-0.123373), (46475,-0.163258), (46476,-0.319272), (46477,-0.315038), (46478,-0.476625), (46479,-0.522553), (46480,-0.698072), (46481,-0.384949), (46482,-0.172151), (46483,-0.220401), (46484,-0.347618), (46485,-0.191025), (46486,-0.247171), (46487,-0.298209), (46488,-0.541085), (46489,-0.235858), (46490,-0.048144), (46491,-0.108004), (46492,-0.278420), (46493,-0.265820), (46494,-0.407432), (46495,-0.485413), (46496,-0.622849), (46497,-0.379393), (46498,-0.111787), (46499,-0.200914), (46500,-0.343922), (46501,-0.254216), (46502,-0.286675), (46503,-0.344218), (46504,-0.642366), (46505,-0.409599), (46506,-0.115981), (46507,-0.254344), (46508,-0.285406), (46509,-0.525026), (46510,-0.492921), (46511,-0.649862), (46512,-0.734812), (46513,-0.490893), (46514,-0.240938), (46515,-0.365832), (46516,-0.439630), (46517,-0.505063), (46518,-0.321069), (46519,-0.470114), (46520,-0.528583), (46521,-0.727334), (46522,-0.047251), (46523,-0.171218), (46524,-0.223646), (46525,-0.393598), (46526,-0.350804), (46527,-0.550945), (46528,-0.588976), (46529,-0.772861), (46530,-0.087213), (46531,-0.227429), (46532,-0.280326), (46533,-0.430304), (46534,-0.206823), (46535,-0.348435), (46536,-0.408765), (46537,-0.616801), (46538,0.074890), (46539,-0.063009), (46540,-0.126588), (46541,-0.263561), (46542,-0.271399), (46543,-0.432059), (46544,-0.490529), (46545,-0.640501), (46546,0.033076), (46547,-0.118292), (46548,-0.173049), (46549,-0.335563), (46550,-0.105119), (46551,-0.286218), (46552,-0.524441), (46553,-0.657231), (46554,0.020058), (46555,-0.149888), (46556,-0.232516), (46557,-0.371341), (46558,-0.368960), (46559,-0.498963), (46560,-0.560220), (46561,-0.712521), (46562,-0.031512), (46563,-0.182880), (46564,-0.232527), (46565,-0.416406), (46566,-0.161341), (46567,-0.344299), (46568,-0.416238), (46569,-0.548095), (46570,0.112933), (46571,-0.028679), (46572,-0.109910), (46573,-0.294259), (46574,-0.290945), (46575,-0.401906), (46576,-0.465022), (46577,-0.574117), (46578,0.085520), (46579,-0.026368), (46580,-0.113172), (46581,-0.245029), (46582,-0.027590), (46583,-0.182672), (46584,-0.394891), (46585,-0.555551), (46586,0.118489), (46587,-0.021734), (46588,-0.096922), (46589,-0.238071), (46590,-0.251019), (46591,-0.382418), (46592,-0.441815), (46593,-0.621517), (46594,0.044627), (46595,-0.078407), (46596,-0.132237), (46597,-0.304970), (46598,-0.070807), (46599,-0.209169), (46600,-0.452046), (46601,-0.586225), (46602,0.068766), (46603,-0.095144), (46604,-0.161040), (46605,-0.283147), (46606,-0.274730), (46607,-0.406593), (46608,-0.487818), (46609,-0.662880), (46610,0.041817), (46611,-0.143922), (46612,-0.179630), (46613,-0.325889), (46614,-0.090799), (46615,-0.264465), (46616,-0.401437), (46617,-0.135684), (46618,-0.290771), (46619,0.059978), (46620,-0.092317), (46621,-0.096905), (46622,-0.248736), (46623,-0.351802), (46624,-0.500847), (46625,-0.202583), (46626,-0.363243), (46627,-0.028286), (46628,-0.164325), (46629,-0.015164), (46630,-0.186507), (46631,-0.160901), (46632,-0.497602), (46633,-0.202595), (46634,0.034818), (46635,0.004683), (46636,-0.147612), (46637,-0.129439), (46638,-0.319360), (46639,-0.362038), (46640,-0.533381), (46641,-0.275066), (46642,-0.013033), (46643,-0.014371), (46644,-0.184781), (46645,-0.009145), (46646,-0.062506), (46647,-0.153956), (46648,-0.520387), (46649,-0.207721), (46650,-0.001899), (46651,-0.065941), (46652,-0.239601), (46653,-0.206569), (46654,-0.392770), (46655,-0.438698), (46656,-0.587280), (46657,-0.305741), (46658,-0.036281), (46659,-0.080812), (46660,-0.266087), (46661,-0.140620), (46662,-0.193980), (46663,-0.232939), (46664,-0.517618), (46665,-0.235616), (46666,0.018059), (46667,-0.050167), (46668,-0.238228), (46669,-0.222378), (46670,-0.392331), (46671,-0.438722), (46672,-0.614241), (46673,-0.331775), (46674,-0.082284), (46675,-0.137967), (46676,-0.303737), (46677,-0.125778), (46678,-0.184248), (46679,-0.273839), (46680,-0.366679), (46681,-0.062842), (46682,-0.216996), (46683,0.143045), (46684,-0.018542), (46685,0.027032), (46686,-0.145701), (46687,-0.210676), (46688,-0.402921), (46689,-0.132527), (46690,-0.282969), (46691,0.067317), (46692,-0.114238), (46693,0.061860), (46694,-0.111342), (46695,-0.112674), (46696,-0.642610), (46697,0.078811), (46698,-0.087885), (46699,-0.163544), (46700,-0.286578), (46701,-0.311604), (46702,-0.464368), (46703,-0.523765), (46704,-0.648195), (46705,-0.001093), (46706,-0.161290), (46707,-0.216504), (46708,-0.368805), (46709,-0.168085), (46710,-0.268822), (46711,-0.318932), (46712,-0.503744), (46713,-0.220808), (46714,0.031464), (46715,-0.024683), (46716,-0.202989), (46717,-0.201077), (46718,-0.389139), (46719,-0.430884), (46720,-0.736934), (46721,-0.476760), (46722,-0.232378), (46723,-0.294097), (46724,-0.429210), (46725,-0.299091), (46726,-0.362207), (46727,-0.382123), (46728,-0.642181), (46729,-0.316980), (46730,-0.099078), (46731,-0.176126), (46732,-0.301947), (46733,-0.301889), (46734,-0.471372), (46735,-0.514513), (46736,-0.676100), (46737,-0.403390), (46738,-0.113949), (46739,-0.159413), (46740,-0.351658), (46741,-0.225721), (46742,-0.285124), (46743,-0.315260), (46744,-0.548844), (46745,-0.677450), (46746,0.020740), (46747,-0.176144), (46748,-0.269917), (46749,-0.424071), (46750,-0.398002), (46751,-0.551693), (46752,-0.627815), (46753,-0.760141), (46754,-0.054048), (46755,-0.189161), (46756,-0.308482), (46757,-0.443595), (46758,-0.244728), (46759,-0.377981), (46760,-0.492193), (46761,-0.644494), (46762,0.016540), (46763,-0.124145), (46764,-0.161707), (46765,-0.346989), (46766,-0.367832), (46767,-0.547997), (46768,-0.560018), (46769,-0.727648), (46770,-0.046639), (46771,-0.178502), (46772,-0.251831), (46773,-0.425960), (46774,-0.171828), (46775,-0.323660), (46776,-0.553061), (46777,-0.679814), (46778,0.012340), (46779,-0.162252), (46780,-0.210503), (46781,-0.363731), (46782,-0.431487), (46783,-0.562417), (46784,-0.625996), (46785,-0.739744), (46786,-0.049449), (46787,-0.202671), (46788,-0.306199), (46789,-0.468250), (46790,-0.263354), (46791,-0.419831), (46792,-0.495483), (46793,-0.677972), (46794,0.016963), (46795,-0.133009), (46796,-0.217490), (46797,-0.399978), (46798,-0.411999), (46799,-0.548971), (46800,-0.592576), (46801,-0.740694), (46802,-0.022059), (46803,-0.212913), (46804,-0.247225), (46805,-0.417178), (46806,-0.168613), (46807,-0.316731), (46808,-0.619989), (46809,-0.734200), (46810,-0.058764), (46811,-0.153464), (46812,-0.258383), (46813,-0.438555), (46814,-0.412022), (46815,-0.581505), (46816,-0.626500), (46817,-0.779264), (46818,-0.074105), (46819,-0.238478), (46820,-0.279766), (46821,-0.465504), (46822,-0.197434), (46823,-0.343693), (46824,-0.455117), (46825,-0.597656), (46826,0.043866), (46827,-0.099143), (46828,-0.141820), (46829,-0.294579), (46830,-0.291271), (46831,-0.451468), (46832,-0.528053), (46833,-0.660373), (46834,0.041531), (46835,-0.139561), (46836,-0.239834), (46837,-0.369373), (46838,-0.138930), (46839,-0.310736), (46840,-0.389174), (46841,-0.530793), (46842,0.119095), (46843,-0.010444), (46844,-0.060085), (46845,-0.228642), (46846,-0.276429), (46847,-0.399463), (46848,-0.453750), (46849,-0.643208), (46850,0.049410), (46851,-0.107068), (46852,-0.160428), (46853,-0.285785), (46854,-0.070670), (46855,-0.220178), (46856,-0.435183), (46857,-0.570759), (46858,0.062404), (46859,-0.074562), (46860,-0.097729), (46861,-0.291833), (46862,-0.342407), (46863,-0.457545), (46864,-0.519264), (46865,-0.665986), (46866,0.012693), (46867,-0.138212), (46868,-0.170670), (46869,-0.349439), (46870,-0.150116), (46871,-0.327032), (46872,-0.449603), (46873,-0.155058), (46874,-0.293884), (46875,0.052689), (46876,-0.085674), (46877,-0.085152), (46878,-0.247203), (46879,-0.347945), (46880,-0.505813), (46881,-0.238212), (46882,-0.335235), (46883,-0.033252), (46884,-0.174870), (46885,-0.000162), (46886,-0.157566), (46887,-0.111529), (46888,-0.536018), (46889,-0.270271), (46890,-0.071875), (46891,-0.116406), (46892,-0.249196), (46893,-0.209658), (46894,-0.395866), (46895,-0.469195), (46896,-0.585729), (46897,-0.300471), (46898,-0.080709), (46899,-0.114558), (46900,-0.252457), (46901,-0.109802), (46902,-0.151084), (46903,-0.245320), (46904,-0.511884), (46905,-0.235455), (46906,0.005678), (46907,-0.037464), (46908,-0.195338), (46909,-0.210608), (46910,-0.381018), (46911,-0.431592), (46912,-0.570424), (46913,-0.322322), (46914,-0.076550), (46915,-0.142916), (46916,-0.296607), (46917,-0.135367), (46918,-0.207312), (46919,-0.255563), (46920,-0.469635), (46921,-0.191346), (46922,0.017270), (46923,-0.034701), (46924,-0.197678), (46925,-0.179505), (46926,-0.362000), (46927,-0.387953), (46928,-0.558362), (46929,-0.273574), (46930,-0.040337), (46931,-0.091374), (46932,-0.268290), (46933,-0.120989), (46934,-0.210579), (46935,-0.226783), (46936,-0.326129), (46937,-0.030651), (46938,-0.201067), (46939,0.130640), (46940,-0.043952), (46941,-0.030425), (46942,-0.185507), (46943,-0.243976), (46944,-0.391631), (46945,-0.096154), (46946,-0.264247), (46947,0.088826), (46948,-0.047214), (46949,0.054102), (46950,-0.140466), (46951,-0.086989), (46952,-0.480822), (46953,-0.193247), (46954,0.062751), (46955,-0.023589), (46956,-0.179604), (46957,-0.161431), (46958,-0.331383), (46959,-0.374988), (46960,-0.521246), (46961,-0.259212), (46962,-0.033415), (46963,-0.103494), (46964,-0.240930), (46965,-0.073190), (46966,-0.154421), (46967,-0.176655), (46968,-0.482705), (46969,-0.230427), (46970,0.005133), (46971,-0.073775), (46972,-0.238149), (46973,-0.188855), (46974,-0.369027), (46975,-0.431673), (46976,-0.832012), (46977,-0.533284), (46978,-0.308414), (46979,-0.356664), (46980,-0.475985), (46981,-0.317532), (46982,-0.404799), (46983,-0.479994), (46984,-0.637398), (46985,-0.374901), (46986,-0.142134), (46987,-0.188062), (46988,-0.357545), (46989,-0.296642), (46990,-0.465662), (46991,-0.542710), (46992,-0.701974), (46993,-0.415325), (46994,-0.176516), (46995,-0.213621), (46996,-0.378458), (46997,-0.236266), (46998,-0.308668), (46999,-0.313256), (47000,-0.584467), (47001,-0.722366), (47002,-0.064582), (47003,-0.178793), (47004,-0.236336), (47005,-0.424861), (47006,-0.448497), (47007,-0.625413), (47008,-0.643006), (47009,-0.788801), (47010,-0.112439), (47011,-0.272630), (47012,-0.303229), (47013,-0.455993), (47014,-0.243664), (47015,-0.362052), (47016,-0.471617), (47017,-0.621126), (47018,0.061737), (47019,-0.086382), (47020,-0.177362), (47021,-0.327803), (47022,-0.354220), (47023,-0.515807), (47024,-0.553838), (47025,-0.724718), (47026,-0.021881), (47027,-0.194151), (47028,-0.226609), (47029,-0.407708), (47030,-0.189800), (47031,-0.345814), (47032,-0.656504), (47033,-0.833883), (47034,-0.154271), (47035,-0.289847), (47036,-0.369218), (47037,-0.481570), (47038,-0.482908), (47039,-0.627307), (47040,-0.715507), (47041,-0.891026), (47042,-0.177970), (47043,-0.350240), (47044,-0.399887), (47045,-0.534530), (47046,-0.314306), (47047,-0.447095), (47048,-0.467939), (47049,-0.621166), (47050,0.047300), (47051,-0.127762), (47052,-0.174153), (47053,-0.365001), (47054,-0.380741), (47055,-0.476368), (47056,-0.547380), (47057,-0.718722), (47058,-0.027495), (47059,-0.155175), (47060,-0.188560), (47061,-0.348757), (47062,-0.110875), (47063,-0.232055), (47064,-0.547855), (47065,-0.715941), (47066,-0.021001), (47067,-0.147291), (47068,-0.236881), (47069,-0.367811), (47070,-0.363107), (47071,-0.553028), (47072,-0.601742), (47073,-0.775871), (47074,-0.116697), (47075,-0.279217), (47076,-0.294951), (47077,-0.465830), (47078,-0.212156), (47079,-0.372816), (47080,-0.418280), (47081,-0.611451), (47082,0.073270), (47083,-0.066488), (47084,-0.121702), (47085,-0.285149), (47086,-0.291597), (47087,-0.478268), (47088,-0.550207), (47089,-0.682997), (47090,-0.027072), (47091,-0.184013), (47092,-0.212289), (47093,-0.346012), (47094,-0.103489), (47095,-0.259497), (47096,-0.245507), (47097,-0.378296), (47098,-0.121842), (47099,0.093280), (47100,0.068253), (47101,-0.112382), (47102,-0.123933), (47103,-0.286453), (47104,-0.606892), (47105,-0.323030), (47106,-0.515738), (47107,-0.123649), (47108,-0.298705), (47109,-0.165342), (47110,-0.318100), (47111,-0.278562), (47112,-0.485672), (47113,-0.660264), (47114,-0.378725), (47115,-0.154318), (47116,-0.196526), (47117,-0.348827), (47118,-0.331117), (47119,-0.526611), (47120,-0.554430), (47121,-0.702079), (47122,-0.462343), (47123,-0.229113), (47124,-0.292692), (47125,-0.431055), (47126,-0.270748), (47127,-0.325962), (47128,-0.569301), (47129,-0.342571), (47130,-0.472574), (47131,-0.122288), (47132,-0.259254), (47133,-0.275458), (47134,-0.444014), (47135,-0.504337), (47136,-0.639913), (47137,-0.376489), (47138,-0.541796), (47139,-0.218911), (47140,-0.360060), (47141,-0.196503), (47142,-0.352518), (47143,-0.338991), (47144,-0.738859), (47145,-0.448034), (47146,-0.237096), (47147,-0.309961), (47148,-0.447860), (47149,-0.448735), (47150,-0.628437), (47151,-0.684121), (47152,-0.799259), (47153,-0.490312), (47154,-0.286343), (47155,-0.361995), (47156,-0.563531), (47157,-0.403225), (47158,-0.428714), (47159,-0.493684), (47160,-0.636692), (47161,-0.311491), (47162,-0.467968), (47163,-0.142303), (47164,-0.302957), (47165,-0.276888), (47166,-0.466346), (47167,-0.524353), (47168,-0.672934), (47169,-0.393249), (47170,-0.535331), (47171,-0.239390), (47172,-0.379612), (47173,-0.233238), (47174,-0.392038), (47175,-0.412882), (47176,-0.628350), (47177,-0.347275), (47178,-0.483314), (47179,-0.172051), (47180,-0.310414), (47181,-0.287131), (47182,-0.440822), (47183,-0.510438), (47184,-0.683171), (47185,-0.406278), (47186,-0.552073), (47187,-0.173916), (47188,-0.298347), (47189,-0.154295), (47190,-0.326101), (47191,-0.297709), (47192,-0.552658), (47193,-0.300849), (47194,-0.452681), (47195,-0.109364), (47196,-0.256549), (47197,-0.237913), (47198,-0.432480), (47199,-0.483054), (47200,-0.644178), (47201,-0.362169), (47202,-0.574388), (47203,-0.219919), (47204,-0.376403), (47205,-0.249070), (47206,-0.405084), (47207,-0.375302), (47208,-0.728259), (47209,-0.414672), (47210,-0.171217), (47211,-0.193920), (47212,-0.376872), (47213,-0.356845), (47214,-0.517969), (47215,-0.566683), (47216,-0.725021), (47217,-0.445335), (47218,-0.194453), (47219,-0.245027), (47220,-0.383390), (47221,-0.237942), (47222,-0.328465), (47223,-0.352095), (47224,-0.784487), (47225,-0.521057), (47226,-0.265529), (47227,-0.311920), (47228,-0.487445), (47229,-0.454407), (47230,-0.645261), (47231,-0.711164), (47232,-1.093850), (47233,-0.418415), (47234,-0.533553), (47235,-0.557189), (47236,-0.712270), (47237,-0.487399), (47238,-0.639230), (47239,-0.735327), (47240,-0.947076), (47241,-0.269323), (47242,-0.417905), (47243,-0.484734), (47244,-0.643998), (47245,-0.703864), (47246,-0.815283), (47247,-0.872826), (47248,-1.065533), (47249,-0.414255), (47250,-0.526143), (47251,-0.566029), (47252,-0.730872), (47253,-0.451650), (47254,-0.604877), (47255,-0.685182), (47256,-0.726000), (47257,-0.918244), (47258,-0.259070), (47259,-0.379781), (47260,-0.405270), (47261,-0.557102), (47262,-0.562623), (47263,-0.743252), (47264,-0.802185), (47265,-0.979564), (47266,-0.248856), (47267,-0.406730), (47268,-0.482852), (47269,-0.632360), (47270,-0.377759), (47271,-0.554674), (47272,-0.888125), (47273,-0.578252), (47274,-0.307859), (47275,-0.444832), (47276,-0.514911), (47277,-0.706691), (47278,-0.682946), (47279,-0.840350), (47280,-0.872809), (47281,-0.666053), (47282,-0.421671), (47283,-0.567929), (47284,-0.587382), (47285,-0.704844), (47286,-0.563579), (47287,-0.705661), (47288,-0.919733), (47289,-0.672101), (47290,-0.403567), (47291,-0.560508), (47292,-0.603650), (47293,-0.775456), (47294,-0.776794), (47295,-0.915157), (47296,-0.979663), (47297,-0.771980), (47298,-0.460247), (47299,-0.638090), (47300,-0.678444), (47301,-0.765248), (47302,-0.646281), (47303,-0.741908), (47304,-0.830108), (47305,-0.580153), (47306,-0.293968), (47307,-0.470414), (47308,-0.537249), (47309,-0.691404), (47310,-0.676944), (47311,-0.831568), (47312,-0.891428), (47313,-0.656338), (47314,-0.379908), (47315,-0.528027), (47316,-0.619940), (47317,-0.678410), (47318,-0.561296), (47319,-0.723347), (47320,-0.786463), (47321,-0.933184), (47322,-0.253572), (47323,-0.425848), (47324,-0.489891), (47325,-0.650545), (47326,-0.670461), (47327,-0.776777), (47328,-0.856148), (47329,-0.965713), (47330,-0.304679), (47331,-0.451401), (47332,-0.510804), (47333,-0.651020), (47334,-0.422899), (47335,-0.541287), (47336,-0.632737), (47337,-0.819408), (47338,-0.161161), (47339,-0.305560), (47340,-0.320830), (47341,-0.498679), (47342,-0.527882), (47343,-0.632337), (47344,-0.687094), (47345,-0.846358), (47346,-0.180678), (47347,-0.324150), (47348,-0.375187), (47349,-0.565108), (47350,-0.356962), (47351,-0.455375), (47352,-0.524991), (47353,-0.669859), (47354,-0.001862), (47355,-0.156017), (47356,-0.255826), (47357,-0.375604), (47358,-0.394131), (47359,-0.537139), (47360,-0.570988), (47361,-0.720966), (47362,-0.067828), (47363,-0.257286), (47364,-0.300891), (47365,-0.422065), (47366,-0.203700), (47367,-0.352745), (47368,-0.597938), (47369,-0.727478), (47370,-0.068303), (47371,-0.220135), (47372,-0.248874), (47373,-0.434619), (47374,-0.453139), (47375,-0.601257), (47376,-0.653228), (47377,-0.832930), (47378,-0.132879), (47379,-0.294466), (47380,-0.341784), (47381,-0.484330), (47382,-0.282683), (47383,-0.437764), (47384,-0.815805), (47385,-0.546808), (47386,-0.268519), (47387,-0.342781), (47388,-0.515520), (47389,-0.527534), (47390,-0.689591), (47391,-0.718330), (47392,-0.859479), (47393,-0.566795), (47394,-0.293145), (47395,-0.382272), (47396,-0.611680), (47397,-0.437434), (47398,-0.501014), (47399,-0.500956), (47400,-0.702029), (47401,-0.438135), (47402,-0.207692), (47403,-0.243400), (47404,-0.387799), (47405,-0.404466), (47406,-0.567449), (47407,-0.629632), (47408,-0.777287), (47409,-0.497602), (47410,-0.230464), (47411,-0.274532), (47412,-0.457021), (47413,-0.274416), (47414,-0.361220), (47415,-0.396929), (47416,-0.681608), (47417,-0.386600), (47418,-0.162656), (47419,-0.234131), (47420,-0.387822), (47421,-0.337602), (47422,-0.534956), (47423,-0.559976), (47424,-0.693235), (47425,-0.420056), (47426,-0.161271), (47427,-0.220668), (47428,-0.418491), (47429,-0.248429), (47430,-0.305039), (47431,-0.344461), (47432,-0.595696), (47433,-0.327626), (47434,-0.070238), (47435,-0.128708), (47436,-0.309807), (47437,-0.295817), (47438,-0.496420), (47439,-0.537238), (47440,-0.698362), (47441,-0.405671), (47442,-0.166404), (47443,-0.195607), (47444,-0.374846), (47445,-0.212679), (47446,-0.283228), (47447,-0.348667), (47448,-0.737390), (47449,-0.427517), (47450,-0.211932), (47451,-0.282481), (47452,-0.458464), (47453,-0.448193), (47454,-0.607457), (47455,-0.664530), (47456,-0.798710), (47457,-0.542255), (47458,-0.293227), (47459,-0.338691), (47460,-0.503998), (47461,-0.308388), (47462,-0.386363), (47463,-0.424394), (47464,-0.819160), (47465,-0.128865), (47466,-0.283483), (47467,-0.366574), (47468,-0.484498), (47469,-0.489550), (47470,-0.652533), (47471,-0.707283), (47472,-0.840073), (47473,-0.152565), (47474,-0.313688), (47475,-0.386091), (47476,-0.525849), (47477,-0.324203), (47478,-0.454670), (47479,-0.489909), (47480,-0.802922), (47481,-0.142821), (47482,-0.326706), (47483,-0.414436), (47484,-0.579737), (47485,-0.588971), (47486,-0.710615), (47487,-0.776981), (47488,-0.926952), (47489,-0.624975), (47490,-0.409397), (47491,-0.453001), (47492,-0.617838), (47493,-0.460318), (47494,-0.495563), (47495,-0.567502), (47496,-0.982705), (47497,-0.304946), (47498,-0.460034), (47499,-0.496206), (47500,-0.679164), (47501,-0.661918), (47502,-0.817005), (47503,-0.877329), (47504,-1.033806), (47505,-0.363023), (47506,-0.482337), (47507,-0.551490), (47508,-0.703791), (47509,-0.472414), (47510,-0.626105), (47511,-0.744029), (47512,-0.845235), (47513,-0.570196), (47514,-0.304449), (47515,-0.373601), (47516,-0.503141), (47517,-0.498437), (47518,-0.701363), (47519,-0.761229), (47520,-0.950218), (47521,-0.663569), (47522,-0.407578), (47523,-0.463724), (47524,-0.628098), (47525,-0.461285), (47526,-0.518365), (47527,-0.567543), (47528,-0.882415), (47529,-0.663117), (47530,-0.347665), (47531,-0.474419), (47532,-0.552394), (47533,-0.732559), (47534,-0.727861), (47535,-0.871796), (47536,-0.948381), (47537,-0.724901), (47538,-0.406668), (47539,-0.567329), (47540,-0.627652), (47541,-0.722815), (47542,-0.576447), (47543,-0.709236), (47544,-0.890329), (47545,-0.596711), (47546,-0.351865), (47547,-0.378751), (47548,-0.535229), (47549,-0.522165), (47550,-0.694435), (47551,-0.729680), (47552,-0.930753), (47553,-0.643172), (47554,-0.371852), (47555,-0.437285), (47556,-0.616993), (47557,-0.474332), (47558,-0.546277), (47559,-0.585235), (47560,-0.827641), (47561,-0.603234), (47562,-0.324018), (47563,-0.438229), (47564,-0.493906), (47565,-0.669895), (47566,-0.650332), (47567,-0.848149), (47568,-0.890358), (47569,-0.637153), (47570,-0.376515), (47571,-0.532993), (47572,-0.585890), (47573,-0.638787), (47574,-0.477083), (47575,-0.643780), (47576,-0.812336), (47577,-0.553089), (47578,-0.338437), (47579,-0.400157), (47580,-0.529233), (47581,-0.497591), (47582,-0.715377), (47583,-0.752482), (47584,-0.903387), (47585,-0.624634), (47586,-0.353314), (47587,-0.415960), (47588,-0.561292), (47589,-0.457190), (47590,-0.529592), (47591,-0.551832), (47592,-0.620521), (47593,-0.692460), (47594,-0.034676), (47595,-0.217170), (47596,-0.262165), (47597,-0.452556), (47598,-0.449242), (47599,-0.605726), (47600,-0.658153), (47601,-0.799302), (47602,-0.135951), (47603,-0.297069), (47604,-0.346252), (47605,-0.515272), (47606,-0.267640), (47607,-0.454775), (47608,-0.651195), (47609,-0.400314), (47610,-0.149895), (47611,-0.168415), (47612,-0.329076), (47613,-0.333201), (47614,-0.526835), (47615,-0.597384), (47616,-0.695797), (47617,-0.411008), (47618,-0.156407), (47619,-0.233918), (47620,-0.353702), (47621,-0.224979), (47622,-0.272767), (47623,-0.319628), (47624,-0.575039), (47625,-0.740346), (47626,-0.075129), (47627,-0.248332), (47628,-0.305869), (47629,-0.458633), (47630,-0.454392), (47631,-0.590438), (47632,-0.656334), (47633,-0.810958), (47634,-0.108585), (47635,-0.282250), (47636,-0.327245), (47637,-0.493015), (47638,-0.266284), (47639,-0.430195), (47640,-0.757603), (47641,-0.524373), (47642,-0.292070), (47643,-0.323132), (47644,-0.435020), (47645,-0.443322), (47646,-0.644858), (47647,-0.692646), (47648,-0.834258), (47649,-0.548536), (47650,-0.344103), (47651,-0.366807), (47652,-0.551155), (47653,-0.404317), (47654,-0.511559), (47655,-0.541695), (47656,-0.682380), (47657,-0.406414), (47658,-0.182933), (47659,-0.213069), (47660,-0.343536), (47661,-0.358343), (47662,-0.514357), (47663,-0.564461), (47664,-0.735804), (47665,-0.447296), (47666,-0.166220), (47667,-0.246525), (47668,-0.437372), (47669,-0.248268), (47670,-0.343895), (47671,-0.387969), (47672,-0.683794), (47673,-0.403182), (47674,-0.109564), (47675,-0.151778), (47676,-0.307786), (47677,-0.270571), (47678,-0.509728), (47679,-0.572844), (47680,-0.696341), (47681,-0.405510), (47682,-0.182962), (47683,-0.226104), (47684,-0.377008), (47685,-0.265937), (47686,-0.305829), (47687,-0.376841), (47688,-0.609028), (47689,-0.371152), (47690,-0.143025), (47691,-0.210787), (47692,-0.364478), (47693,-0.346305), (47694,-0.495350), (47695,-0.598415), (47696,-0.740954), (47697,-0.444550), (47698,-0.156975), (47699,-0.245169), (47700,-0.392360), (47701,-0.219042), (47702,-0.331857), (47703,-0.358743), (47704,-0.703340), (47705,-0.429233), (47706,-0.168596), (47707,-0.208487), (47708,-0.384470), (47709,-0.365370), (47710,-0.588272), (47711,-0.634199), (47712,-0.761879), (47713,-0.468725), (47714,-0.266615), (47715,-0.338091), (47716,-0.490849), (47717,-0.356553), (47718,-0.366714), (47719,-0.458627), (47720,-0.792542), (47721,-0.127795), (47722,-0.291242), (47723,-0.374796), (47724,-0.501080), (47725,-0.522386), (47726,-0.671901), (47727,-0.748949), (47728,-0.888238), (47729,-0.183548), (47730,-0.328874), (47731,-0.375734), (47732,-0.534998), (47733,-0.318023), (47734,-0.467995), (47735,-0.532971), (47736,-0.728928), (47737,-0.476650), (47738,-0.237384), (47739,-0.272622), (47740,-0.449538), (47741,-0.406750), (47742,-0.617110), (47743,-0.676976), (47744,-1.138622), (47745,-0.472479), (47746,-0.589477), (47747,-0.666988), (47748,-0.806747), (47749,-0.574907), (47750,-0.730921), (47751,-0.769416), (47752,-0.834392), (47753,-0.619270), (47754,-0.318220), (47755,-0.487240), (47756,-0.533167), (47757,-0.718912), (47758,-0.738366), (47759,-0.912958), (47760,-0.870164), (47761,-0.656909), (47762,-0.393015), (47763,-0.515586), (47764,-0.563373), (47765,-0.619056), (47766,-0.452244), (47767,-0.611508), (47768,-0.867853), (47769,-0.608612), (47770,-0.335895), (47771,-0.498872), (47772,-0.555489), (47773,-0.752373), (47774,-0.723054), (47775,-0.887891), (47776,-0.943574), (47777,-0.651353), (47778,-0.373527), (47779,-0.558802), (47780,-0.633997), (47781,-0.669242), (47782,-0.527514), (47783,-0.679809), (47784,-0.777295), (47785,-0.552887), (47786,-0.303402), (47787,-0.445478), (47788,-0.502551), (47789,-0.686899), (47790,-0.656654), (47791,-0.811272), (47792,-0.895289), (47793,-0.621646), (47794,-0.318736), (47795,-0.475683), (47796,-0.509996), (47797,-0.557320), (47798,-0.383074), (47799,-0.535375), (47800,-0.864644), (47801,-0.640700), (47802,-0.375879), (47803,-0.561161), (47804,-0.581541), (47805,-0.766352), (47806,-0.737497), (47807,-0.865640), (47808,-0.924110), (47809,-0.709452), (47810,-0.433023), (47811,-0.630840), (47812,-0.681877), (47813,-0.762645), (47814,-0.576327), (47815,-0.711903), (47816,-0.716028), (47817,-0.453067), (47818,-0.207288), (47819,-0.373522), (47820,-0.394365), (47821,-0.617267), (47822,-0.582838), (47823,-0.756504), (47824,-0.797322), (47825,-0.551080), (47826,-0.283480), (47827,-0.419519), (47828,-0.467770), (47829,-0.503479), (47830,-0.379865), (47831,-0.528447), (47832,-0.861898), (47833,-0.603584), (47834,-0.305320), (47835,-0.446005), (47836,-0.502615), (47837,-0.678135), (47838,-0.662285), (47839,-0.809940), (47840,-0.919505), (47841,-0.673263), (47842,-0.389864), (47843,-0.529623), (47844,-0.594129), (47845,-0.686506), (47846,-0.538278), (47847,-0.696615), (47848,-0.766231), (47849,-0.492124), (47850,-0.229164), (47851,-0.377276), (47852,-0.457117), (47853,-0.638209), (47854,-0.604244), (47855,-0.772800), (47856,-0.837306), (47857,-0.594320), (47858,-0.273302), (47859,-0.445571), (47860,-0.535161), (47861,-0.596881), (47862,-0.442147), (47863,-0.599088), (47864,-0.574879), (47865,-0.762013), (47866,-0.038738), (47867,-0.195216), (47868,-0.240680), (47869,-0.405987), (47870,-0.453768), (47871,-0.584698), (47872,-0.658966), (47873,-0.763885), (47874,-0.120033), (47875,-0.255146), (47876,-0.316865), (47877,-0.469630), (47878,-0.217815), (47879,-0.376615), (47880,-0.609273), (47881,-0.723014), (47882,-0.035969), (47883,-0.197563), (47884,-0.255563), (47885,-0.443161), (47886,-0.396660), (47887,-0.566606), (47888,-0.631112), (47889,-0.758329), (47890,-0.100082), (47891,-0.245877), (47892,-0.318279), (47893,-0.442246), (47894,-0.237343), (47895,-0.394291), (47896,-0.658062), (47897,-0.368164), (47898,-0.123781), (47899,-0.186897), (47900,-0.358240), (47901,-0.347500), (47902,-0.547640), (47903,-0.555478), (47904,-0.742613), (47905,-0.493584), (47906,-0.273823), (47907,-0.309531), (47908,-0.438608), (47909,-0.294093), (47910,-0.336771), (47911,-0.412886), (47912,-0.841095), (47913,-0.183781), (47914,-0.290553), (47915,-0.332304), (47916,-0.505037), (47917,-0.542142), (47918,-0.674469), (47919,-0.715750), (47920,-0.843894), (47921,-0.181470), (47922,-0.317039), (47923,-0.384802), (47924,-0.530597), (47925,-0.290861), (47926,-0.464526), (47927,-0.504412), (47928,-0.636275), (47929,-0.324542), (47930,-0.130791), (47931,-0.171146), (47932,-0.361067), (47933,-0.344284), (47934,-0.504018), (47935,-0.579207), (47936,-0.736147), (47937,-0.441603), (47938,-0.182825), (47939,-0.232929), (47940,-0.393590), (47941,-0.250471), (47942,-0.327983), (47943,-0.378093), (47944,-0.640938), (47945,-0.358472), (47946,-0.114090), (47947,-0.206467), (47948,-0.355975), (47949,-0.351741), (47950,-0.541198), (47951,-0.574121), (47952,-0.730598), (47953,-0.477393), (47954,-0.222792), (47955,-0.271506), (47956,-0.403363), (47957,-0.278359), (47958,-0.356341), (47959,-0.386940), (47960,-0.614481), (47961,-0.328296), (47962,-0.115504), (47963,-0.165144), (47964,-0.323482), (47965,-0.338752), (47966,-0.493840), (47967,-0.536048), (47968,-0.689739), (47969,-0.417029), (47970,-0.162891), (47971,-0.211605), (47972,-0.387131), (47973,-0.216599), (47974,-0.311305), (47975,-0.373025), (47976,-0.744559), (47977,-0.058447), (47978,-0.219571), (47979,-0.263176), (47980,-0.389459), (47981,-0.397297), (47982,-0.520801), (47983,-0.566729), (47984,-0.746894), (47985,-0.089580), (47986,-0.268818), (47987,-0.369091), (47988,-0.509777), (47989,-0.231488), (47990,-0.376813), (47991,-0.439002), (47992,-0.886253), (47993,-0.229865), (47994,-0.359869), (47995,-0.448526), (47996,-0.598504), (47997,-0.611451), (47998,-0.730309), (47999,-0.811533), (48000,-0.844456), (48001,-0.986074), (48002,-0.335723), (48003,-0.487554), (48004,-0.526982), (48005,-0.685783), (48006,-0.450223), (48007,-0.621566), (48008,-0.765038), (48009,-0.888072), (48010,-0.227971), (48011,-0.377479), (48012,-0.444315), (48013,-0.582208), (48014,-0.595162), (48015,-0.740487), (48016,-0.768300), (48017,-0.952648), (48018,-0.317631), (48019,-0.469463), (48020,-0.565089), (48021,-0.677904), (48022,-0.427022), (48023,-0.581640), (48024,-0.726509), (48025,-0.798447), (48026,-0.507153), (48027,-0.254874), (48028,-0.399273), (48029,-0.454493), (48030,-0.662993), (48031,-0.618809), (48032,-0.805943), (48033,-0.839335), (48034,-0.594490), (48035,-0.271605), (48036,-0.443881), (48037,-0.513496), (48038,-0.590544), (48039,-0.434421), (48040,-0.878885), (48041,-0.525806), (48042,-0.679967), (48043,-0.396099), (48044,-0.526102), (48045,-0.571103), (48046,-0.757311), (48047,-0.750747), (48048,-0.897005), (48049,-0.563444), (48050,-0.733391), (48051,-0.450455), (48052,-0.558630), (48053,-0.533025), (48054,-0.750353), (48055,-0.601192), (48056,-0.806442), (48057,-0.841224), (48058,-0.620993), (48059,-0.346423), (48060,-0.491749), (48061,-0.520494), (48062,-0.726671), (48063,-0.709894), (48064,-0.873804), (48065,-0.915549), (48066,-0.638656), (48067,-0.360831), (48068,-0.513125), (48069,-0.582747), (48070,-0.605914), (48071,-0.510171), (48072,-0.657826), (48073,-0.724655), (48074,-0.505821), (48075,-0.209880), (48076,-0.385869), (48077,-0.478709), (48078,-0.616145), (48079,-0.592399), (48080,-0.776277), (48081,-0.805486), (48082,-0.596871), (48083,-0.360848), (48084,-0.492711), (48085,-0.532139), (48086,-0.608717), (48087,-0.431229), (48088,-0.761887), (48089,-0.800852), (48090,-0.573195), (48091,-0.318130), (48092,-0.462992), (48093,-0.485232), (48094,-0.667257), (48095,-0.647224), (48096,-0.799525), (48097,-0.879360), (48098,-0.655416), (48099,-0.412430), (48100,-0.564261), (48101,-0.574422), (48102,-0.668196), (48103,-0.509285), (48104,-0.704779), (48105,-0.737238), (48106,-0.492856), (48107,-0.197378), (48108,-0.347356), (48109,-0.377955), (48110,-0.592491), (48111,-0.583610), (48112,-0.716863), (48113,-0.797168), (48114,-0.558358), (48115,-0.252198), (48116,-0.420755), (48117,-0.451817), (48118,-0.540944), (48119,-0.412221), (48120,-0.702010), (48121,-0.721463), (48122,-0.486373), (48123,-0.196469), (48124,-0.328332), (48125,-0.370077), (48126,-0.560461), (48127,-0.543221), (48128,-0.696449), (48129,-0.728908), (48130,-0.486379), (48131,-0.206236), (48132,-0.381292), (48133,-0.461597), (48134,-0.485226), (48135,-0.323987), (48136,-0.670443), (48137,-0.703366), (48138,-0.491964), (48139,-0.249441), (48140,-0.391986), (48141,-0.426768), (48142,-0.610647), (48143,-0.586438), (48144,-0.751744), (48145,-0.792099), (48146,-0.575587), (48147,-0.235051), (48148,-0.428228), (48149,-0.471833), (48150,-0.549808), (48151,-0.405299), (48152,-0.580355), (48153,-0.717321), (48154,-0.452038), (48155,-0.235063), (48156,-0.273558), (48157,-0.427719), (48158,-0.416978), (48159,-0.589248), (48160,-0.656077), (48161,-0.832529), (48162,-0.496175), (48163,-0.262482), (48164,-0.339067), (48165,-0.482539), (48166,-0.335701), (48167,-0.409499), (48168,-0.647260), (48169,-0.780513), (48170,-0.113906), (48171,-0.258311), (48172,-0.295410), (48173,-0.453747), (48174,-0.508034), (48175,-0.674267), (48176,-0.715085), (48177,-0.887824), (48178,-0.202639), (48179,-0.313131), (48180,-0.375314), (48181,-0.561522), (48182,-0.345937), (48183,-0.471294), (48184,-0.726243), (48185,-0.864605), (48186,-0.156196), (48187,-0.334508), (48188,-0.405983), (48189,-0.554101), (48190,-0.580517), (48191,-0.750934), (48192,-0.760631), (48193,-0.904567), (48194,-0.229131), (48195,-0.376322), (48196,-0.427823), (48197,-0.570368), (48198,-0.304151), (48199,-0.432295), (48200,-0.620826), (48201,-0.757329), (48202,-0.056815), (48203,-0.226298), (48204,-0.277335), (48205,-0.470513), (48206,-0.503898), (48207,-0.658979), (48208,-0.717449), (48209,-0.929668), (48210,-0.239373), (48211,-0.342896), (48212,-0.406475), (48213,-0.554593), (48214,-0.319967), (48215,-0.460189), (48216,-0.436907), (48217,-0.615212), (48218,-0.339246), (48219,-0.118095), (48220,-0.189100), (48221,-0.336755), (48222,-0.306510), (48223,-0.527088), (48224,-0.563724), (48225,-0.686294), (48226,-0.387103), (48227,-0.128789), (48228,-0.222556), (48229,-0.368351), (48230,-0.247061), (48231,-0.358486), (48232,-0.724447), (48233,-0.509796), (48234,-0.248695), (48235,-0.358723), (48236,-0.413937), (48237,-0.536507), (48238,-0.523914), (48239,-0.712438), (48240,-0.775554), (48241,-0.539531), (48242,-0.241737), (48243,-0.408897), (48244,-0.438570), (48245,-0.520264), (48246,-0.361347), (48247,-0.537336), (48248,-0.656187), (48249,-0.784794), (48250,-0.120980), (48251,-0.294176), (48252,-0.359615), (48253,-0.494258), (48254,-0.514638), (48255,-0.641855), (48256,-0.897737), (48257,-1.054214), (48258,-0.414082), (48259,-0.522251), (48260,-0.594659), (48261,-0.705614), (48262,-0.500718), (48263,-0.645117), (48264,-0.822496), (48265,-0.986406), (48266,-0.269174), (48267,-0.393598), (48268,-0.481798), (48269,-0.641062), (48270,-0.629395), (48271,-0.784939), (48272,-0.840623), (48273,-1.012429), (48274,-0.349541), (48275,-0.539926), (48276,-0.603969), (48277,-0.696809), (48278,-0.452426), (48279,-0.614947), (48280,-0.910771), (48281,-0.954839), (48282,-0.734615), (48283,-0.449356), (48284,-0.583079), (48285,-0.649908), (48286,-0.828214), (48287,-0.825369), (48288,-0.953513), (48289,-0.982258), (48290,-0.734163), (48291,-0.462837), (48292,-0.625820), (48293,-0.727489), (48294,-0.778990), (48295,-0.606604), (48296,-0.970249), (48297,-0.616244), (48298,-0.761113), (48299,-0.502328), (48300,-0.632795), (48301,-0.734001), (48302,-0.871437), (48303,-0.880201), (48304,-1.033892), (48305,-0.671997), (48306,-0.811287), (48307,-0.559008), (48308,-0.677396), (48309,-0.703355), (48310,-0.811061), (48311,-0.691630), (48312,-0.846248), (48313,-0.874061), (48314,-0.637574), (48315,-0.376474), (48316,-0.507867), (48317,-0.562624), (48318,-0.747898), (48319,-0.751090), (48320,-0.879703), (48321,-0.939100), (48322,-0.718406), (48323,-0.418752), (48324,-0.578949), (48325,-0.626266), (48326,-0.732582), (48327,-0.569952), (48328,-0.762196), (48329,-0.820666), (48330,-0.571638), (48331,-0.289635), (48332,-0.441003), (48333,-0.471602), (48334,-0.681962), (48335,-0.691196), (48336,-0.817943), (48337,-0.870377), (48338,-0.616702), (48339,-0.359321), (48340,-0.497683), (48341,-0.546861), (48342,-0.613226), (48343,-0.481254), (48344,-0.895988), (48345,-0.943775), (48346,-0.692893), (48347,-0.396489), (48348,-0.570618), (48349,-0.629551), (48350,-0.804607), (48351,-0.760887), (48352,-0.923870), (48353,-0.985590), (48354,-0.731452), (48355,-0.468491), (48356,-0.670491), (48357,-0.701554), (48358,-0.773962), (48359,-0.620155), (48360,-0.778492), (48361,-0.830456), (48362,-0.617201), (48363,-0.347271), (48364,-0.484243), (48365,-0.547816), (48366,-0.732165), (48367,-0.713528), (48368,-0.876512), (48369,-0.899678), (48370,-0.679917), (48371,-0.373757), (48372,-0.552532), (48373,-0.626794), (48374,-0.651820), (48375,-0.531457), (48376,-0.698153), (48377,-0.757556), (48378,-0.510851), (48379,-0.266932), (48380,-0.401118), (48381,-0.447509), (48382,-0.643466), (48383,-0.651311), (48384,-0.732072), (48385,-0.853716), (48386,-0.604688), (48387,-0.320825), (48388,-0.505174), (48389,-0.558071), (48390,-0.634656), (48391,-0.469703), (48392,-0.769241), (48393,-0.845362), (48394,-0.571719), (48395,-0.311545), (48396,-0.459200), (48397,-0.534852), (48398,-0.700158), (48399,-0.677339), (48400,-0.860760), (48401,-0.949418), (48402,-0.691567), (48403,-0.394236), (48404,-0.581834), (48405,-0.618006), (48406,-0.660684), (48407,-0.504560), (48408,-0.620624), (48409,-0.771066), (48410,-0.531793), (48411,-0.276265), (48412,-0.312900), (48413,-0.480993), (48414,-0.458638), (48415,-0.615585), (48416,-0.664762), (48417,-0.852824), (48418,-0.567102), (48419,-0.345951), (48420,-0.360288), (48421,-0.508870), (48422,-0.342527), (48423,-0.422361), (48424,-0.752099), (48425,-0.903931), (48426,-0.254512), (48427,-0.378009), (48428,-0.419754), (48429,-0.584598), (48430,-0.599405), (48431,-0.760059), (48432,-0.819925), (48433,-0.979189), (48434,-0.320478), (48435,-0.445835), (48436,-0.529389), (48437,-0.706768), (48438,-0.469819), (48439,-0.594712), (48440,-0.776274), (48441,-0.905808), (48442,-0.297729), (48443,-0.449097), (48444,-0.489915), (48445,-0.607839), (48446,-0.646334), (48447,-0.808391), (48448,-0.850136), (48449,-0.996858), (48450,-0.334897), (48451,-0.463974), (48452,-0.540559), (48453,-0.734656), (48454,-0.451257), (48455,-0.566859), (48456,-0.697795), (48457,-0.868668), (48458,-0.192775), (48459,-0.359935), (48460,-0.366846), (48461,-0.560017), (48462,-0.577611), (48463,-0.746631), (48464,-0.794418), (48465,-0.930921), (48466,-0.248986), (48467,-0.415219), (48468,-0.496913), (48469,-0.638062), (48470,-0.406222), (48471,-0.546444), (48472,-0.592835), (48473,-0.774860), (48474,-0.505864), (48475,-0.245689), (48476,-0.317628), (48477,-0.425797), (48478,-0.396941), (48479,-0.606837), (48480,-0.662057), (48481,-0.831077), (48482,-0.533276), (48483,-0.225727), (48484,-0.305561), (48485,-0.447173), (48486,-0.290586), (48487,-0.327222), (48488,-0.800953), (48489,-0.522194), (48490,-0.258307), (48491,-0.417107), (48492,-0.450030), (48493,-0.620439), (48494,-0.650112), (48495,-0.775006), (48496,-0.858560), (48497,-0.633689), (48498,-0.337278), (48499,-0.516517), (48500,-0.522965), (48501,-0.618128), (48502,-0.399294), (48503,-0.579002), (48504,-0.657440), (48505,-0.801845), (48506,-0.156603), (48507,-0.261522), (48508,-0.366904), (48509,-0.502017), (48510,-0.494990), (48511,-0.677485), (48512,-0.957048), (48513,-1.087984), (48514,-0.421841), (48515,-0.571349), (48516,-0.649330), (48517,-0.775151), (48518,-0.547024), (48519,-0.708611), (48520,-0.870667), (48521,-1.009493), (48522,-0.344277), (48523,-0.498901), (48524,-0.560157), (48525,-0.685514), (48526,-0.703571), (48527,-0.875840), (48528,-0.956608), (48529,-1.096830), (48530,-0.420005), (48531,-0.575086), (48532,-0.674895), (48533,-0.807221), (48534,-0.570735), (48535,-0.718390), (48536,-0.722045), (48537,-0.781911), (48538,-0.925847), (48539,-0.276428), (48540,-0.434296), (48541,-0.498338), (48542,-0.631591), (48543,-0.616211), (48544,-0.753641), (48545,-0.846951), (48546,-0.989026), (48547,-0.305237), (48548,-0.420839), (48549,-0.513215), (48550,-0.647865), (48551,-0.447609), (48552,-0.810784), (48553,-0.879936), (48554,-0.615586), (48555,-0.329400), (48556,-0.492378), (48557,-0.579181), (48558,-0.724513), (48559,-0.684975), (48560,-0.826124), (48561,-0.884131), (48562,-0.627670), (48563,-0.351704), (48564,-0.518400), (48565,-0.553646), (48566,-0.647419), (48567,-0.443449), (48568,-0.831709), (48569,-0.921299), (48570,-0.711294), (48571,-0.418603), (48572,-0.537454), (48573,-0.650738), (48574,-0.806753), (48575,-0.796012), (48576,-0.945984), (48577,-1.036037), (48578,-0.780046), (48579,-0.481782), (48580,-0.637796), (48581,-0.694406), (48582,-0.783533), (48583,-0.633909), (48584,-0.818721), (48585,-0.864648), (48586,-0.584506), (48587,-0.320612), (48588,-0.472450), (48589,-0.515591), (48590,-0.702726), (48591,-0.671547), (48592,-0.820129), (48593,-0.861874), (48594,-0.604023), (48595,-0.316911), (48596,-0.484071), (48597,-0.579697), (48598,-0.672544), (48599,-0.514090), (48600,-0.669178), (48601,-0.718355), (48602,-0.875760), (48603,-0.224018), (48604,-0.368423), (48605,-0.434789), (48606,-0.597303), (48607,-0.591208), (48608,-0.781593), (48609,-0.825661), (48610,-0.945445), (48611,-0.299276), (48612,-0.430676), (48613,-0.502151), (48614,-0.638191), (48615,-0.458836), (48616,-0.634362), (48617,-0.677503), (48618,-0.785208), (48619,-0.124638), (48620,-0.281578), (48621,-0.368382), (48622,-0.483520), (48623,-0.469993), (48624,-0.608819), (48625,-0.690050), (48626,-0.836309), (48627,-0.135795), (48628,-0.274158), (48629,-0.334951), (48630,-0.441729), (48631,-0.250765), (48632,-0.467161), (48633,-0.530277), (48634,-0.702546), (48635,-0.013642), (48636,-0.171516), (48637,-0.230912), (48638,-0.400395), (48639,-0.450042), (48640,-0.591191), (48641,-0.650124), (48642,-0.784774), (48643,-0.118167), (48644,-0.255133), (48645,-0.346583), (48646,-0.504457), (48647,-0.242887), (48648,-0.569832), (48649,-0.633411), (48650,-0.756915), (48651,-0.093094), (48652,-0.209159), (48653,-0.274598), (48654,-0.416211), (48655,-0.422658), (48656,-0.575886), (48657,-0.614845), (48658,-0.802443), (48659,-0.172529), (48660,-0.301142), (48661,-0.330808), (48662,-0.510511), (48663,-0.300968), (48664,-0.648352), (48665,-0.811798), (48666,-0.533973), (48667,-0.288664), (48668,-0.348530), (48669,-0.502221), (48670,-0.483585), (48671,-0.670256), (48672,-0.733829), (48673,-0.866619), (48674,-0.602268), (48675,-0.339307), (48676,-0.408460), (48677,-0.578869), (48678,-0.442720), (48679,-0.482605), (48680,-0.543862), (48681,-0.671542), (48682,-0.468036), (48683,-0.219014), (48684,-0.278874), (48685,-0.402841), (48686,-0.392100), (48687,-0.576912), (48688,-0.626089), (48689,-0.763525), (48690,-0.493132), (48691,-0.249676), (48692,-0.291427), (48693,-0.441399), (48694,-0.314999), (48695,-0.359537), (48696,-0.531343), (48697,-0.674352), (48698,-0.416037), (48699,-0.186984), (48700,-0.268678), (48701,-0.399608), (48702,-0.369819), (48703,-0.552778), (48704,-0.610314), (48705,-0.760756), (48706,-0.474107), (48707,-0.193032), (48708,-0.247782), (48709,-0.442349), (48710,-0.313626), (48711,-0.359091), (48712,-0.513245), (48713,-0.639535), (48714,-0.380288), (48715,-0.154490), (48716,-0.238501), (48717,-0.342494), (48718,-0.368916), (48719,-0.501700), (48720,-0.603832), (48721,-0.742664), (48722,-0.474594), (48723,-0.273411), (48724,-0.307724), (48725,-0.483712), (48726,-0.333625), (48727,-0.396271), (48728,-0.626142), (48729,-0.783083), (48730,-0.483429), (48731,-0.226504), (48732,-0.319814), (48733,-0.449811), (48734,-0.453936), (48735,-0.607627), (48736,-0.632653), (48737,-0.796100), (48738,-0.508055), (48739,-0.278075), (48740,-0.356519), (48741,-0.501845), (48742,-0.374518), (48743,-0.422306), (48744,-0.593648), (48745,-0.773350), (48746,-0.062618), (48747,-0.220485), (48748,-0.276632), (48749,-0.468413), (48750,-0.447917), (48751,-0.600218), (48752,-0.650792), (48753,-0.825384), (48754,-0.109072), (48755,-0.223747), (48756,-0.289649), (48757,-0.474924), (48758,-0.242621), (48759,-0.393989), (48760,-0.735799), (48761,-0.877881), (48762,-0.189910), (48763,-0.348241), (48764,-0.413680), (48765,-0.565048), (48766,-0.554307), (48767,-0.705212), (48768,-0.788766), (48769,-0.800317), (48770,-0.588452), (48771,-0.291584), (48772,-0.477323), (48773,-0.566450), (48774,-0.634675), (48775,-0.464149), (48776,-0.719098), (48777,-0.734368), (48778,-0.529936), (48779,-0.241891), (48780,-0.394192), (48781,-0.425718), (48782,-0.627254), (48783,-0.627660), (48784,-0.781351), (48785,-0.823565), (48786,-0.601481), (48787,-0.319942), (48788,-0.506607), (48789,-0.572973), (48790,-0.604041), (48791,-0.496683), (48792,-0.803660), (48793,-0.861197), (48794,-0.593590), (48795,-0.351068), (48796,-0.454597), (48797,-0.528858), (48798,-0.704847), (48799,-0.678778), (48800,-0.864980), (48801,-0.910444), (48802,-0.705085), (48803,-0.425399), (48804,-0.563762), (48805,-0.649639), (48806,-0.719718), (48807,-0.558485), (48808,-0.774417), (48809,-0.543967), (48810,-0.558774), (48811,-0.724544), (48812,-0.427213), (48813,-0.619457), (48814,-0.664452), (48815,-0.827435), (48816,-0.778605), (48817,-0.556521), (48818,-0.559249), (48819,-0.703654), (48820,-0.479247), (48821,-0.548399), (48822,-0.634270), (48823,-0.778675), (48824,-0.736344), (48825,-0.876103), (48826,-0.498410), (48827,-0.638632), (48828,-0.343624), (48829,-0.498242), (48830,-0.594802), (48831,-0.745706), (48832,-0.731246), (48833,-0.864963), (48834,-0.517933), (48835,-0.677197), (48836,-0.371500), (48837,-0.535411), (48838,-0.508415), (48839,-0.662569), (48840,-0.590515), (48841,-0.725164), (48842,-0.388347), (48843,-0.551330), (48844,-0.277218), (48845,-0.389569), (48846,-0.520969), (48847,-0.677910), (48848,-0.672742), (48849,-0.820860), (48850,-0.482184), (48851,-0.655386), (48852,-0.347366), (48853,-0.483876), (48854,-0.455947), (48855,-0.607315), (48856,-0.697368), (48857,-0.873821), (48858,-0.516102), (48859,-0.686982), (48860,-0.422625), (48861,-0.527544), (48862,-0.636645), (48863,-0.799629), (48864,-0.777736), (48865,-0.956975), (48866,-0.627127), (48867,-0.774319), (48868,-0.525754), (48869,-0.677585), (48870,-0.633871), (48871,-0.783842), (48872,-0.630042), (48873,-0.785123), (48874,-0.434373), (48875,-0.558804), (48876,-0.316745), (48877,-0.454637), (48878,-0.516827), (48879,-0.663085), (48880,-0.655131), (48881,-0.809749), (48882,-0.487334), (48883,-0.654494), (48884,-0.372955), (48885,-0.515037), (48886,-0.458311), (48887,-0.620361), (48888,-0.532051), (48889,-0.646726), (48890,-0.270892), (48891,-0.450131), (48892,-0.172305), (48893,-0.321813), (48894,-0.404904), (48895,-0.581356), (48896,-0.591517), (48897,-0.763787), (48898,-0.428366), (48899,-0.541644), (48900,-0.277757), (48901,-0.426339), (48902,-0.416525), (48903,-0.559997), (48904,-0.558549), (48905,-0.682510), (48906,-0.342443), (48907,-0.492421), (48908,-0.200193), (48909,-0.385005), (48910,-0.456950), (48911,-0.629219), (48912,-0.652386), (48913,-0.801430), (48914,-0.401446), (48915,-0.556527), (48916,-0.349308), (48917,-0.491383), (48918,-0.462528), (48919,-0.604610), (48920,-0.552993), (48921,-0.590098), (48922,-0.731711), (48923,-0.036770), (48924,-0.199753), (48925,-0.253577), (48926,-0.393793), (48927,-0.449476), (48928,-0.578553), (48929,-0.571525), (48930,-0.766093), (48931,-0.084157), (48932,-0.251787), (48933,-0.273094), (48934,-0.442577), (48935,-0.209347), (48936,-0.655201), (48937,-0.723427), (48938,-0.484617), (48939,-0.223516), (48940,-0.356306), (48941,-0.412453), (48942,-0.592155), (48943,-0.580488), (48944,-0.741142), (48945,-0.770814), (48946,-0.548730), (48947,-0.252325), (48948,-0.407413), (48949,-0.470059), (48950,-0.551290), (48951,-0.383088), (48952,-0.620848), (48953,-0.687683), (48954,-0.419144), (48955,-0.134355), (48956,-0.300125), (48957,-0.358125), (48958,-0.525291), (48959,-0.489466), (48960,-0.651053), (48961,-0.748540), (48962,-0.559436), (48963,-0.295079), (48964,-0.427868), (48965,-0.450571), (48966,-0.527156), (48967,-0.374746), (48968,-0.647346), (48969,-0.763410), (48970,-0.458184), (48971,-0.172925), (48972,-0.329872), (48973,-0.392519), (48974,-0.566648), (48975,-0.559157), (48976,-0.733286), (48977,-0.814981), (48978,-0.529729), (48979,-0.215210), (48980,-0.372150), (48981,-0.433870), (48982,-0.482121), (48983,-0.371976), (48984,-0.448098), (48985,-0.482880), (48986,-0.646790), (48987,-0.018273), (48988,-0.151989), (48989,-0.169120), (48990,-0.338603), (48991,-0.397999), (48992,-0.505704), (48993,-0.607837), (48994,-0.743876), (48995,-0.100031), (48996,-0.237003), (48997,-0.307546), (48998,-0.454737), (48999,-0.205709), (49000,-0.771405), (49001,-0.381176), (49002,-0.516289), (49003,-0.288625), (49004,-0.433030), (49005,-0.537949), (49006,-0.678165), (49007,-0.648383), (49008,-0.752839), (49009,-0.417881), (49010,-0.596187), (49011,-0.308612), (49012,-0.462766), (49013,-0.446916), (49014,-0.609430), (49015,-0.489073), (49016,-0.684567), (49017,-0.691941), (49018,-0.461961), (49019,-0.168807), (49020,-0.322961), (49021,-0.349384), (49022,-0.553700), (49023,-0.509053), (49024,-0.516897), (49025,-0.207018), (49026,-0.334698), (49027,-0.041544), (49028,-0.177589), (49029,-0.137119), (49030,-0.339582), (49031,-0.232224), (49032,-0.442120), (49033,-0.062573), (49034,-0.239489), (49035,0.019289), (49036,-0.169699), (49037,-0.219809), (49038,-0.371641), (49039,-0.345108), (49040,-0.461173), (49041,-0.152696), (49042,-0.291986), (49043,-0.011837), (49044,-0.175747), (49045,-0.154324), (49046,-0.288973), (49047,-0.142599), (49048,-0.398017), (49049,-0.184292), (49050,-0.239975), (49051,-0.360686), (49052,-0.085184), (49053,-0.271385), (49054,-0.327069), (49055,-0.512350), (49056,-0.470489), (49057,-0.188480), (49058,-0.271101), (49059,-0.412257), (49060,-0.125602), (49061,-0.220771), (49062,-0.293637), (49063,-0.406915), (49064,-0.281912), (49065,-0.054254), (49066,-0.084390), (49067,-0.248300), (49068,0.015593), (49069,-0.156676), (49070,-0.232798), (49071,-0.387885), (49072,-0.395260), (49073,-0.156450), (49074,-0.236285), (49075,-0.328662), (49076,-0.059202), (49077,-0.126031), (49078,-0.182177), (49079,-0.344228), (49080,-0.305623), (49081,-0.075636), (49082,-0.168946), (49083,-0.320314), (49084,-0.029020), (49085,-0.201289), (49086,-0.248150), (49087,-0.419956), (49088,-0.406892), (49089,-0.145785), (49090,-0.167098), (49091,-0.318930), (49092,-0.038317), (49093,-0.106080), (49094,-0.158507), (49095,-0.331709), (49096,-0.258728), (49097,0.007952), (49098,-0.055164), (49099,-0.203745), (49100,0.055965), (49101,-0.097262), (49102,-0.129721), (49103,-0.298741), (49104,-0.271275), (49105,-0.022253), (49106,-0.113234), (49107,-0.244170), (49108,0.002072), (49109,-0.089841), (49110,-0.138556), (49111,-0.255553), (49112,-0.344680), (49113,-0.112377), (49114,-0.168060), (49115,-0.320355), (49116,-0.030450), (49117,-0.192044), (49118,-0.268159), (49119,-0.439038), (49120,-0.422262), (49121,-0.196921), (49122,-0.280475), (49123,-0.444849), (49124,-0.146585), (49125,-0.197622), (49126,-0.226831), (49127,-0.396778), (49128,-0.247623), (49129,-0.049226), (49130,-0.097477), (49131,-0.254881), (49132,0.022011), (49133,-0.154435), (49134,-0.222660), (49135,-0.399112), (49136,-0.398128), (49137,-0.153282), (49138,-0.209429), (49139,-0.344072), (49140,-0.055564), (49141,-0.143764), (49142,-0.196198), (49143,-0.368467), (49144,-0.092501), (49145,-0.274056), (49146,0.094345), (49147,-0.075608), (49148,0.205004), (49149,0.046667), (49150,-0.046173), (49151,-0.194292), (49152,-0.111554), (49153,-0.318194), (49154,0.069712), (49155,-0.082120), (49156,0.173408), (49157,-0.001184), (49158,0.044396), (49159,-0.111618), (49160,-0.170551), (49161,-0.311706), (49162,0.067847), (49163,-0.089094), (49164,0.163178), (49165,0.035967), (49166,-0.043404), (49167,-0.211497), (49168,-0.227231), (49169,-0.345155), (49170,-0.005558), (49171,-0.173182), (49172,0.085133), (49173,-0.040224), (49174,-0.032270), (49175,-0.173419), (49176,-0.232816), (49177,-0.225795), (49178,-0.027398), (49179,0.216057), (49180,0.084194), (49181,0.080070), (49182,-0.146082), (49183,-0.154383), (49184,-0.291355), (49185,-0.336350), (49186,-0.100797), (49187,0.185852), (49188,-0.004069), (49189,-0.038382), (49190,-0.117290), (49191,0.036975), (49192,-0.398197), (49193,-0.056271), (49194,-0.184878), (49195,0.077613), (49196,-0.082114), (49197,-0.139188), (49198,-0.274764), (49199,-0.260773), (49200,-0.374052), (49201,-0.029808), (49202,-0.217406), (49203,0.062743), (49204,-0.055182), (49205,-0.022150), (49206,-0.178158), (49207,-0.039222), (49208,-0.176188), (49209,-0.257883), (49210,-0.001891), (49211,0.301482), (49212,0.092050), (49213,0.057737), (49214,-0.118715), (49215,-0.107511), (49216,-0.271885), (49217,-0.315026), (49218,-0.097588), (49219,0.184421), (49220,0.012615), (49221,-0.024954), (49222,-0.105721), (49223,0.077347), (49224,-0.205009), (49225,-0.279271), (49226,-0.018634), (49227,0.266162), (49228,0.124080), (49229,0.060500), (49230,-0.121525), (49231,-0.148405), (49232,-0.282591), (49233,-0.346633), (49234,-0.102251), (49235,0.163496), (49236,0.013055), (49237,-0.009649), (49238,-0.062076), (49239,0.053172), (49240,-0.201777), (49241,-0.236559), (49242,0.003641), (49243,0.328379), (49244,0.129172), (49245,0.087421), (49246,-0.110860), (49247,-0.122881), (49248,-0.256134), (49249,-0.328072), (49250,-0.027022), (49251,0.192739), (49252,0.033939), (49253,-0.008739), (49254,-0.126663), (49255,0.078239), (49256,-0.286802), (49257,0.017034), (49258,-0.164521), (49259,0.110049), (49260,-0.021808), (49261,-0.076565), (49262,-0.241865), (49263,-0.195364), (49264,-0.329080), (49265,0.010060), (49266,-0.112974), (49267,0.147200), (49268,0.011160), (49269,0.009822), (49270,-0.093237), (49271,0.017364), (49272,-0.265918), (49273,0.079258), (49274,-0.090688), (49275,0.187601), (49276,0.039019), (49277,-0.107702), (49278,-0.287411), (49279,-0.233008), (49280,-0.486560), (49281,-0.250080), (49282,-0.114851), (49283,-0.269939), (49284,-0.339091), (49285,-0.407780), (49286,-0.116485), (49287,-0.286432), (49288,-0.446629), (49289,-0.099592), (49290,-0.250960), (49291,-0.255549), (49292,-0.401344), (49293,-0.480252), (49294,-0.593530), (49295,-0.342185), (49296,-0.455463), (49297,-0.104714), (49298,-0.267691), (49299,-0.099025), (49300,-0.280123), (49301,-0.280992), (49302,-0.400313), (49303,-0.146175), (49304,-0.297079), (49305,-0.386670), (49306,-0.155293), (49307,-0.108786), (49308,-0.285702), (49309,-0.351604), (49310,-0.537349), (49311,-0.228402), (49312,-0.413214), (49313,-0.458215), (49314,-0.212900), (49315,-0.054916), (49316,-0.181669), (49317,-0.223878), (49318,-0.306968), (49319,-0.026356), (49320,-0.358874), (49321,-0.010912), (49322,-0.163213), (49323,-0.147363), (49324,-0.295481), (49325,-0.399003), (49326,-0.523897), (49327,-0.254900), (49328,-0.352850), (49329,0.002546), (49330,-0.173907), (49331,-0.029855), (49332,-0.151963), (49333,-0.128680), (49334,-0.267506), (49335,-0.050531), (49336,-0.423925), (49337,-0.088505), (49338,-0.240799), (49339,-0.254680), (49340,-0.427413), (49341,-0.531405), (49342,-0.668841), (49343,-0.390088), (49344,-0.550279), (49345,-0.199993), (49346,-0.341605), (49347,-0.166440), (49348,-0.298296), (49349,-0.332615), (49350,-0.433814), (49351,-0.171317), (49352,-0.394682), (49353,-0.088059), (49354,-0.188338), (49355,-0.162732), (49356,-0.342434), (49357,-0.422269), (49358,-0.569460), (49359,-0.299067), (49360,-0.442076), (49361,-0.120587), (49362,-0.276601), (49363,-0.137196), (49364,-0.323861), (49365,-0.292219), (49366,-0.441271), (49367,-0.182486), (49368,-0.340824), (49369,-0.396044), (49370,-0.171636), (49371,-0.164146), (49372,-0.304831), (49373,-0.368874), (49374,-0.532321), (49375,-0.237770), (49376,-0.372419), (49377,-0.412311), (49378,-0.179538), (49379,-0.059644), (49380,-0.230053), (49381,-0.260189), (49382,-0.311226), (49383,-0.037583), (49384,-0.188025), (49385,-0.216301), (49386,-0.018837), (49387,-0.020639), (49388,-0.192445), (49389,-0.242086), (49390,-0.390668), (49391,-0.071966), (49392,-0.244705), (49393,-0.284590), (49394,-0.058792), (49395,0.104301), (49396,-0.053567), (49397,-0.101818), (49398,-0.175153), (49399,0.088271), (49400,-0.164354), (49401,-0.211215), (49402,0.028991), (49403,0.052267), (49404,-0.088882), (49405,-0.137596), (49406,-0.348419), (49407,-0.108219), (49408,-0.133709), (49409,-0.210294), (49410,0.051271), (49411,0.180927), (49412,0.018406), (49413,-0.056319), (49414,-0.119435), (49415,0.128197), (49416,-0.151836), (49417,-0.191257), (49418,0.031754), (49419,0.024379), (49420,-0.099118), (49421,-0.148765), (49422,-0.335900), (49423,-0.035776), (49424,-0.172749), (49425,-0.219140), (49426,-0.001702), (49427,0.106583), (49428,-0.041065), (49429,-0.097212), (49430,-0.202131), (49431,0.128643), (49432,-0.143030), (49433,-0.293935), (49434,0.093978), (49435,-0.039739), (49436,-0.094495), (49437,-0.247254), (49438,-0.008451), (49439,-0.132411), (49440,-0.217362), (49441,-0.353864), (49442,0.157603), (49443,0.032246), (49444,-0.012291), (49445,-0.151581), (49446,0.144823), (49447,-0.005618), (49448,-0.142121), (49449,-0.310214), (49450,0.125544), (49451,-0.047658), (49452,-0.070361), (49453,-0.267252), (49454,-0.002432), (49455,-0.144044), (49456,-0.210873), (49457,-0.371070), (49458,0.177091), (49459,0.022937), (49460,-0.047149), (49461,-0.178542), (49462,0.170817), (49463,0.034778), (49464,-0.159326), (49465,-0.313950), (49466,0.105546), (49467,-0.041176), (49468,-0.098249), (49469,-0.248227), (49470,0.010557), (49471,-0.169152), (49472,-0.199751), (49473,-0.309310), (49474,0.223053), (49475,0.008518), (49476,-0.018832), (49477,-0.175773), (49478,0.123418), (49479,0.033828), (49480,-0.099425), (49481,-0.246154), (49482,0.188671), (49483,0.026621), (49484,-0.056470), (49485,-0.211088), (49486,0.047227), (49487,-0.124580), (49488,-0.160288), (49489,-0.347886), (49490,0.205384), (49491,0.055406), (49492,0.033173), (49493,-0.114945), (49494,0.184245), (49495,0.037523), (49496,-0.115241), (49497,-0.248494), (49498,0.148241), (49499,0.013128), (49500,-0.036976), (49501,-0.172089), (49502,0.090872), (49503,-0.077221), (49504,-0.149623), (49505,-0.293095), (49506,0.243451), (49507,0.063285), (49508,0.037332), (49509,-0.106140), (49510,0.263651), (49511,0.121575), (49512,-0.146848), (49513,0.184859), (49514,0.048356), (49515,0.045622), (49516,-0.097850), (49517,-0.194873), (49518,-0.343918), (49519,-0.099073), (49520,-0.243008), (49521,0.146294), (49522,-0.014829), (49523,0.139904), (49524,0.019194), (49525,0.023434), (49526,-0.126543), (49527,0.174044), (49528,-0.226295), (49529,0.020874), (49530,0.050656), (49531,-0.136479), (49532,-0.228856), (49533,-0.389046), (49534,-0.123299), (49535,-0.271881), (49536,-0.433468), (49537,-0.121272), (49538,-0.255458), (49539,-0.083536), (49540,-0.248372), (49541,-0.223236), (49542,-0.408975), (49543,-0.147410), (49544,-0.405145), (49545,-0.053470), (49546,-0.230385), (49547,-0.209889), (49548,-0.352434), (49549,-0.410898), (49550,-0.614294), (49551,-0.354120), (49552,-0.479477), (49553,-0.153342), (49554,-0.295888), (49555,-0.129538), (49556,-0.252109), (49557,-0.265526), (49558,-0.392737), (49559,-0.106088), (49560,-0.130188), (49561,-0.302457), (49562,0.059908), (49563,-0.074742), (49564,-0.082580), (49565,-0.229771), (49566,-0.335154), (49567,-0.454005), (49568,-0.175715), (49569,-0.356814), (49570,-0.034399), (49571,-0.141641), (49572,-0.028246), (49573,-0.171719), (49574,-0.121029), (49575,-0.288658), (49576,-0.227286), (49577,0.042644), (49578,-0.015363), (49579,-0.152329), (49580,-0.128119), (49581,-0.334302), (49582,-0.382553), (49583,-0.583620), (49584,-0.319263), (49585,-0.040510), (49586,-0.106876), (49587,-0.232696), (49588,-0.106303), (49589,-0.136432), (49590,-0.180043), (49591,-0.336051), (49592,-0.323921), (49593,-0.111122), (49594,-0.155660), (49595,-0.337222), (49596,-0.314403), (49597,-0.467167), (49598,-0.521917), (49599,-0.690010), (49600,-0.380601), (49601,-0.136218), (49602,-0.216516), (49603,-0.383213), (49604,-0.259136), (49605,-0.273943), (49606,-0.333346), (49607,-0.500506), (49608,-0.258911), (49609,-0.044722), (49610,-0.091583), (49611,-0.229476), (49612,-0.208516), (49613,-0.380322), (49614,-0.421147), (49615,-0.630573), (49616,-0.316980), (49617,-0.105585), (49618,-0.127818), (49619,-0.316813), (49620,-0.153720), (49621,-0.245633), (49622,-0.289701), (49623,-0.399729), (49624,-0.140952), (49625,-0.302539), (49626,0.029632), (49627,-0.116163), (49628,-0.107282), (49629,-0.252144), (49630,-0.316187), (49631,-0.497286), (49632,-0.201808), (49633,-0.346213), (49634,-0.008463), (49635,-0.173770), (49636,-0.005104), (49637,-0.182019), (49638,-0.158737), (49639,-0.306385), (49640,-0.062473), (49641,-0.186897), (49642,0.181968), (49643,0.002729), (49644,0.009750), (49645,-0.167629), (49646,-0.249787), (49647,-0.389539), (49648,-0.115896), (49649,-0.268661), (49650,0.075589), (49651,-0.078566), (49652,0.049224), (49653,-0.105857), (49654,-0.081184), (49655,-0.216297), (49656,0.004397), (49657,-0.131179), (49658,0.225143), (49659,0.099786), (49660,0.099844), (49661,-0.061743), (49662,-0.143900), (49663,-0.307347), (49664,-0.043923), (49665,-0.209223), (49666,0.127124), (49667,-0.018671), (49668,0.135599), (49669,-0.028774), (49670,0.017733), (49671,-0.122953), (49672,-0.015131), (49673,-0.194370), (49674,0.149410), (49675,0.050064), (49676,0.016215), (49677,-0.129580), (49678,-0.221957), (49679,-0.369142), (49680,-0.080640), (49681,-0.219929), (49682,0.095053), (49683,-0.019152), (49684,0.174135), (49685,-0.008823), (49686,-0.018521), (49687,-0.146664), (49688,-0.208384), (49689,-0.287755), (49690,-0.015972), (49691,-0.022877), (49692,-0.179360), (49693,-0.213673), (49694,-0.409630), (49695,-0.082105), (49696,-0.257631), (49697,-0.280334), (49698,-0.059640), (49699,0.093234), (49700,-0.057670), (49701,-0.157480), (49702,-0.194585), (49703,0.090210), (49704,-0.088102), (49705,-0.131243), (49706,0.061581), (49707,0.063498), (49708,-0.091589), (49709,-0.071556), (49710,-0.247082), (49711,0.004733), (49712,-0.166146), (49713,-0.193496), (49714,0.025802), (49715,0.182396), (49716,-0.004276), (49717,-0.036728), (49718,-0.101704), (49719,0.191451), (49720,-0.076040), (49721,-0.168423), (49722,0.055521), (49723,0.085773), (49724,-0.048413), (49725,-0.128248), (49726,-0.334888), (49727,0.011215), (49728,-0.221442), (49729,-0.268759), (49730,-0.034133), (49731,0.152648), (49732,-0.008939), (49733,-0.040465), (49734,-0.116586), (49735,0.159843), (49736,-0.085819), (49737,-0.150325), (49738,0.096843), (49739,0.122449), (49740,-0.073515), (49741,-0.123156), (49742,-0.264774), (49743,0.020484), (49744,-0.142963), (49745,-0.174488), (49746,0.019725), (49747,0.193037), (49748,0.021231), (49749,-0.011228), (49750,-0.089666), (49751,0.207202), (49752,-0.177345), (49753,-0.254393), (49754,-0.016047), (49755,-0.000667), (49756,-0.172009), (49757,-0.187280), (49758,-0.350720), (49759,-0.058499), (49760,-0.242384), (49761,-0.314786), (49762,-0.043003), (49763,0.102445), (49764,-0.039637), (49765,-0.130154), (49766,-0.191410), (49767,0.086879), (49768,-0.198733), (49769,0.178960), (49770,0.025269), (49771,0.018821), (49772,-0.130687), (49773,-0.181261), (49774,-0.304295), (49775,-0.065949), (49776,-0.212214), (49777,0.087447), (49778,-0.064385), (49779,0.095922), (49780,-0.056379), (49781,-0.003836), (49782,-0.193287), (49783,0.125409), (49784,-0.300477), (49785,0.030303), (49786,-0.105273), (49787,-0.111721), (49788,-0.242651), (49789,-0.335954), (49790,-0.484072), (49791,-0.236440), (49792,-0.330677), (49793,-0.377068), (49794,-0.169849), (49795,0.003464), (49796,-0.131649), (49797,-0.189649), (49798,-0.247656), (49799,0.010195), (49800,-0.147679), (49801,-0.292077), (49802,0.074464), (49803,-0.070398), (49804,-0.075450), (49805,-0.223568), (49806,-0.289934), (49807,-0.442698), (49808,-0.187634), (49809,-0.325533), (49810,0.000139), (49811,-0.141480), (49812,-0.009971), (49813,-0.152979), (49814,-0.157098), (49815,-0.313575), (49816,-0.136087), (49817,-0.271663), (49818,0.050759), (49819,-0.123370), (49820,-0.101948), (49821,-0.252389), (49822,-0.335943), (49823,-0.446898), (49824,-0.169072), (49825,-0.343665), (49826,0.001048), (49827,-0.136851), (49828,-0.001165), (49829,-0.149284), (49830,-0.151549), (49831,-0.275509), (49832,-0.275915), (49833,-0.040361), (49834,-0.078393), (49835,-0.231621), (49836,-0.220417), (49837,-0.410338), (49838,-0.474844), (49839,-0.625286), (49840,-0.357679), (49841,-0.146277), (49842,-0.195924), (49843,-0.324067), (49844,-0.199521), (49845,-0.251955), (49846,-0.306705), (49847,-0.497559), (49848,-0.237385), (49849,-0.361815), (49850,-0.000377), (49851,-0.134563), (49852,-0.137755), (49853,-0.294696), (49854,-0.384286), (49855,-0.517076), (49856,-0.272694), (49857,-0.422208), (49858,-0.066350), (49859,-0.196816), (49860,-0.024431), (49861,-0.212492), (49862,-0.182246), (49863,-0.363802), (49864,-0.147290), (49865,-0.300518), (49866,0.055804), (49867,-0.096027), (49868,-0.089933), (49869,-0.267312), (49870,-0.335538), (49871,-0.480870), (49872,-0.200721), (49873,-0.367417), (49874,-0.052435), (49875,-0.169896), (49876,-0.056965), (49877,-0.253855), (49878,-0.213384), (49879,-0.321553), (49880,-0.161246), (49881,-0.294036), (49882,0.043245), (49883,-0.106733), (49884,-0.088560), (49885,-0.243641), (49886,-0.305831), (49887,-0.461382), (49888,-0.231395), (49889,-0.376263), (49890,-0.013435), (49891,-0.176419), (49892,-0.057452), (49893,-0.198131), (49894,-0.200402), (49895,-0.356880), (49896,-0.085090), (49897,-0.214630), (49898,0.125437), (49899,-0.018499), (49900,-0.034696), (49901,-0.131719), (49902,-0.225955), (49903,-0.399621), (49904,-0.139447), (49905,-0.272237), (49906,0.052038), (49907,-0.101653), (49908,0.016851), (49909,-0.115939), (49910,-0.079187), (49911,-0.182710), (49912,-0.097186), (49913,-0.255523), (49914,0.089190), (49915,-0.098409), (49916,-0.088138), (49917,-0.244152), (49918,-0.321200), (49919,-0.475818), (49920,-0.094412), (49921,-0.241597), (49922,0.081745), (49923,-0.071019), (49924,0.028906), (49925,-0.087622), (49926,-0.068522), (49927,-0.199922), (49928,-0.051224), (49929,-0.180764), (49930,0.194143), (49931,0.031159), (49932,0.011243), (49933,-0.155454), (49934,-0.233429), (49935,-0.416850), (49936,-0.144134), (49937,-0.310367), (49938,0.047351), (49939,-0.115626), (49940,0.036315), (49941,-0.148960), (49942,-0.082941), (49943,-0.226413), (49944,-0.172943), (49945,-0.277862), (49946,-0.049735), (49947,-0.008807), (49948,-0.154602), (49949,-0.214462), (49950,-0.374190), (49951,-0.112625), (49952,-0.247268), (49953,-0.360083), (49954,-0.123603), (49955,0.053892), (49956,-0.099799), (49957,-0.148977), (49958,-0.180046), (49959,0.098243), (49960,-0.080526), (49961,-0.089297), (49962,0.121179), (49963,0.156997), (49964,-0.027814), (49965,-0.078388), (49966,-0.228823), (49967,0.058752), (49968,-0.113054), (49969,-0.171987), (49970,0.027336), (49971,0.196472), (49972,0.059969), (49973,0.025650), (49974,-0.063940), (49975,0.209703), (49976,-0.162765), (49977,-0.237490), (49978,0.028720), (49979,0.031102), (49980,-0.118407), (49981,-0.140647), (49982,-0.331031), (49983,-0.080613), (49984,-0.229194), (49985,-0.306712), (49986,-0.075335), (49987,0.106336), (49988,-0.025057), (49989,-0.069588), (49990,-0.153142), (49991,0.140939), (49992,-0.137698), (49993,-0.231008), (49994,0.018947), (49995,0.052449), (49996,-0.073371), (49997,-0.106763), (49998,-0.295288), (49999,-0.031864), (50000,-0.217602), (50001,-0.240775), (50002,-0.047018), (50003,0.075662), (50004,-0.070597), (50005,-0.084477), (50006,-0.142947), (50007,0.134416), (50008,-0.127502), (50009,-0.211520), (50010,0.031466), (50011,0.035244), (50012,-0.113808), (50013,-0.134651), (50014,-0.331542), (50015,-0.071367), (50016,-0.224125), (50017,-0.247762), (50018,0.017522), (50019,0.120234), (50020,0.012992), (50021,-0.028290), (50022,-0.139251), (50023,0.142294), (50024,-0.121947), (50025,0.098741), (50026,0.045381), (50027,-0.105054), (50028,-0.136123), (50029,-0.305606), (50030,-0.360819), (50031,-0.562819), (50032,-0.262239), (50033,-0.003455), (50034,-0.071680), (50035,-0.215616), (50036,-0.047876), (50037,-0.098913), (50038,-0.144841), (50039,-0.324080), (50040,-0.186534), (50041,-0.185550), (50042,0.023529), (50043,0.057031), (50044,-0.110592), (50045,-0.196006), (50046,-0.352947), (50047,-0.045860), (50048,-0.319851), (50049,-0.476335), (50050,-0.157633), (50051,-0.311787), (50052,-0.158450), (50053,-0.283807), (50054,-0.283285), (50055,-0.408642), (50056,-0.167510), (50057,-0.304476), (50058,0.020262), (50059,-0.130179), (50060,-0.092038), (50061,-0.236436), (50062,-0.329740), (50063,-0.479254), (50064,-0.182387), (50065,-0.347687), (50066,-0.003907), (50067,-0.135764), (50068,-0.006577), (50069,-0.160269), (50070,-0.139309), (50071,-0.271635), (50072,-0.188898), (50073,-0.360241), (50074,-0.009955), (50075,-0.135775), (50076,-0.105060), (50077,-0.281513), (50078,-0.370176), (50079,-0.500173), (50080,-0.209811), (50081,-0.341668), (50082,-0.048983), (50083,-0.177590), (50084,-0.030289), (50085,-0.191413), (50086,-0.161624), (50087,-0.328784), (50088,-0.090908), (50089,-0.214875), (50090,0.096858), (50091,-0.033139), (50092,-0.067457), (50093,-0.194204), (50094,-0.277295), (50095,-0.415194), (50096,-0.174525), (50097,-0.339368), (50098,-0.024849), (50099,-0.143700), (50100,-0.016374), (50101,-0.116183), (50102,-0.090578), (50103,-0.255414), (50104,-0.240961), (50105,-0.443424), (50106,-0.098248), (50107,-0.261695), (50108,-0.256064), (50109,-0.409291), (50110,-0.489589), (50111,-0.610300), (50112,-0.315756), (50113,-0.479666), (50114,-0.147958), (50115,-0.257060), (50116,-0.132050), (50117,-0.292711), (50118,-0.260136), (50119,-0.450063), (50120,-0.085839), (50121,-0.198190), (50122,0.110293), (50123,-0.032253), (50124,-0.012220), (50125,-0.138047), (50126,-0.264794), (50127,-0.397120), (50128,-0.130903), (50129,-0.274375), (50130,0.045253), (50131,-0.127023), (50132,0.019815), (50133,-0.140839), (50134,-0.127312), (50135,-0.267997), (50136,-0.251221), (50137,-0.362639), (50138,-0.006780), (50139,-0.156295), (50140,-0.157164), (50141,-0.306678), (50142,-0.342387), (50143,-0.544850), (50144,-0.260982), (50145,-0.411423), (50146,-0.032803), (50147,-0.172562), (50148,-0.046162), (50149,-0.228651), (50150,-0.250427), (50151,-0.395753), (50152,-0.413346), (50153,-0.134131), (50154,0.091204), (50155,0.003473), (50156,-0.185521), (50157,-0.170598), (50158,-0.343801), (50159,-0.397624), (50160,-0.543419), (50161,-0.290678), (50162,-0.039326), (50163,-0.080608), (50164,-0.212007), (50165,-0.057737), (50166,-0.138035), (50167,-0.195578), (50168,0.076675), (50169,-0.083522), (50170,-0.112262), (50171,0.118182), (50172,0.097339), (50173,-0.079114), (50174,-0.101353), (50175,-0.267587), (50176,0.056225), (50177,-0.083064), (50178,-0.163369), (50179,0.022486), (50180,0.176293), (50181,0.011450), (50182,-0.009857), (50183,-0.090625), (50184,-0.297728), (50185,-0.031517), (50186,-0.203324), (50187,0.166937), (50188,0.026252), (50189,0.039315), (50190,-0.099047), (50191,-0.198394), (50192,-0.291703), (50193,-0.080765), (50194,-0.220054), (50195,0.136732), (50196,-0.034148), (50197,0.108977), (50198,-0.041001), (50199,-0.014932), (50200,-0.051104), (50201,-0.088672), (50202,-0.236791), (50203,0.184565), (50204,0.016009), (50205,-0.059643), (50206,-0.214267), (50207,0.062162), (50208,-0.077590), (50209,-0.140243), (50210,-0.283715), (50211,0.270952), (50212,0.114938), (50213,0.081552), (50214,-0.070285), (50215,0.211723), (50216,-0.099893), (50217,-0.264273), (50218,0.053039), (50219,-0.082537), (50220,-0.033244), (50221,-0.178576), (50222,-0.249588), (50223,-0.416748), (50224,-0.079004), (50225,-0.239201), (50226,0.069746), (50227,-0.066294), (50228,0.056393), (50229,-0.133528), (50230,-0.076339), (50231,-0.179404), (50232,-0.001909), (50233,-0.035295), (50234,-0.147183), (50235,0.235156), (50236,0.094934), (50237,0.016490), (50238,-0.142774), (50239,0.103931), (50240,-0.049760), (50241,-0.129132), (50242,-0.268890), (50243,0.268588), (50244,0.113037), (50245,0.047605), (50246,-0.092618), (50247,0.267424), (50248,0.094221), (50249,-0.051574), (50250,-0.064521), (50251,0.187294), (50252,0.170163), (50253,0.021118), (50254,-0.092166), (50255,-0.241211), (50256,-0.003798), (50257,-0.152843), (50258,-0.161614), (50259,0.100883), (50260,0.227746), (50261,0.125151), (50262,0.045779), (50263,-0.042415), (50264,0.050542), (50265,0.002754), (50266,-0.163479), (50267,0.238829), (50268,0.084211), (50269,0.025278), (50270,-0.101476), (50271,0.121072), (50272,-0.040045), (50273,-0.071114), (50274,-0.248493), (50275,0.297345), (50276,0.144117), (50277,0.097726), (50278,-0.081513), (50279,0.252055), (50280,0.018934), (50281,-0.127324), (50282,0.214596), (50283,0.041863), (50284,0.080938), (50285,-0.112697), (50286,-0.151198), (50287,-0.269123), (50288,-0.005229), (50289,-0.180291), (50290,0.154666), (50291,0.059040), (50292,0.161288), (50293,0.025242), (50294,0.029947), (50295,-0.087051), (50296,-0.088383), (50297,-0.272268), (50298,0.069189), (50299,-0.122586), (50300,-0.109522), (50301,-0.245098), (50302,-0.332835), (50303,-0.455869), (50304,-0.291843), (50305,-0.440888), (50306,-0.077596), (50307,-0.250799), (50308,-0.127186), (50309,-0.280877), (50310,-0.270136), (50311,-0.410358), (50312,-0.210566), (50313,-0.375409), (50314,-0.024660), (50315,-0.204825), (50316,-0.195944), (50317,-0.342203), (50318,-0.427147), (50319,-0.540425), (50320,-0.268172), (50321,-0.396785), (50322,-0.057645), (50323,-0.239207), (50324,-0.104448), (50325,-0.239554), (50326,-0.250648), (50327,-0.420595), (50328,-0.199437), (50329,-0.327117), (50330,0.000871), (50331,-0.100335), (50332,-0.103527), (50333,-0.253505), (50334,-0.324510), (50335,-0.493530), (50336,-0.229643), (50337,-0.381474), (50338,-0.086930), (50339,-0.206250), (50340,-0.056156), (50341,-0.231682), (50342,-0.207936), (50343,-0.355121), (50344,-0.431706), (50345,-0.143667), (50346,0.091892), (50347,0.054324), (50348,-0.102617), (50349,-0.076085), (50350,-0.256250), (50351,-0.326336), (50352,-0.491636), (50353,-0.229138), (50354,0.018494), (50355,-0.033477), (50356,-0.207143), (50357,-0.066341), (50358,-0.129457), (50359,-0.180957), (50360,-0.634245), (50361,-0.311366), (50362,-0.089282), (50363,-0.128710), (50364,-0.269395), (50365,-0.241467), (50366,-0.419309), (50367,-0.458737), (50368,-0.612428), (50369,-0.330889), (50370,-0.091616), (50371,-0.157519), (50372,-0.314923), (50373,-0.169012), (50374,-0.273468), (50375,-0.357022), (50376,-0.519535), (50377,-0.232887), (50378,0.030074), (50379,-0.037225), (50380,-0.176978), (50381,-0.181566), (50382,-0.384493), (50383,-0.402549), (50384,-0.537662), (50385,-0.255660), (50386,-0.011741), (50387,-0.095295), (50388,-0.242017), (50389,-0.079850), (50390,-0.170837), (50391,-0.225588), (50392,-0.539534), (50393,-0.211539), (50394,-0.007570), (50395,-0.072082), (50396,-0.209975), (50397,-0.214563), (50398,-0.390089), (50399,-0.451345), (50400,-0.598067), (50401,-0.308632), (50402,-0.089798), (50403,-0.178925), (50404,-0.307531), (50405,-0.160693), (50406,-0.227059), (50407,-0.273920), (50408,-0.414606), (50409,-0.092184), (50410,0.134077), (50411,0.103941), (50412,-0.080871), (50413,-0.058051), (50414,-0.267484), (50415,-0.329204), (50416,-0.470816), (50417,-0.202746), (50418,0.034204), (50419,-0.015443), (50420,-0.178884), (50421,-0.077568), (50422,-0.149977), (50423,-0.169424), (50424,-0.199559), (50425,0.077333), (50426,-0.061956), (50427,0.277178), (50428,0.107232), (50429,0.136087), (50430,-0.079382), (50431,-0.156893), (50432,-0.292469), (50433,0.002539), (50434,-0.159512), (50435,0.157794), (50436,0.025937), (50437,0.186244), (50438,0.021401), (50439,0.060475), (50440,-0.233953), (50441,0.044336), (50442,-0.106569), (50443,0.239534), (50444,0.077021), (50445,0.084975), (50446,-0.040382), (50447,-0.176422), (50448,-0.293883), (50449,-0.037892), (50450,-0.192973), (50451,0.136875), (50452,0.010585), (50453,0.181574), (50454,0.003732), (50455,0.020978), (50456,0.106965), (50457,-0.052299), (50458,-0.080581), (50459,0.153119), (50460,0.170828), (50461,-0.007947), (50462,-0.052948), (50463,-0.204779), (50464,0.033567), (50465,-0.129417), (50466,-0.173955), (50467,0.070428), (50468,0.239100), (50469,0.085872), (50470,0.073852), (50471,-0.024098), (50472,0.009397), (50473,-0.154043), (50474,0.162799), (50475,0.002602), (50476,-0.008022), (50477,-0.135702), (50478,-0.244341), (50479,-0.395709), (50480,-0.069574), (50481,-0.234411), (50482,0.070352), (50483,-0.057328), (50484,0.102979), (50485,-0.053035), (50486,-0.030679), (50487,-0.171828), (50488,0.116210), (50489,-0.093679), (50490,-0.138217), (50491,0.112665), (50492,0.140594), (50493,-0.009848), (50494,-0.056702), (50495,-0.267525), (50496,0.076255), (50497,-0.102520), (50498,-0.147978), (50499,0.065277), (50500,0.226054), (50501,0.086758), (50502,0.006924), (50503,-0.095209), (50504,0.128272), (50505,-0.050040), (50506,-0.030007), (50507,0.212979), (50508,0.203281), (50509,-0.001042), (50510,-0.040464), (50511,-0.181613), (50512,0.107359), (50513,-0.112293), (50514,-0.165653), (50515,0.077333), (50516,0.206519), (50517,0.040755), (50518,0.004114), (50519,-0.031595), (50520,0.122212), (50521,-0.017547), (50522,-0.024458), (50523,0.211102), (50524,0.173997), (50525,0.024952), (50526,-0.011690), (50527,-0.179313), (50528,0.113841), (50529,-0.051466), (50530,-0.125727), (50531,0.109363), (50532,0.277572), (50533,0.084394), (50534,0.052405), (50535,-0.038118), (50536,0.046942), (50537,-0.119291), (50538,0.226349), (50539,0.068481), (50540,0.055064), (50541,-0.104664), (50542,-0.117611), (50543,-0.271302), (50544,-0.046431), (50545,-0.187580), (50546,0.156669), (50547,-0.001668), (50548,0.140061), (50549,0.027246), (50550,0.023121), (50551,-0.097127), (50552,-0.092429), (50553,-0.253083), (50554,0.099990), (50555,-0.038836), (50556,-0.048534), (50557,-0.222200), (50558,-0.281596), (50559,-0.433897), (50560,-0.259189), (50561,-0.396161), (50562,-0.071886), (50563,-0.204206), (50564,-0.064338), (50565,-0.168793), (50566,-0.169199), (50567,-0.309884), (50568,-0.070618), (50569,-0.188073), (50570,0.160817), (50571,-0.004490), (50572,-0.003498), (50573,-0.131642), (50574,-0.213336), (50575,-0.397685), (50576,-0.142620), (50577,-0.268910), (50578,0.084162), (50579,-0.115978), (50580,0.072200), (50581,-0.094027), (50582,-0.070751), (50583,-0.214223), (50584,-0.461739), (50585,-0.195529), (50586,0.052567), (50587,-0.003580), (50588,-0.161448), (50589,-0.129806), (50590,-0.334129), (50591,-0.382380), (50592,-0.529565), (50593,-0.214119), (50594,0.028867), (50595,-0.018914), (50596,-0.228810), (50597,-0.102874), (50598,-0.120937), (50599,-0.182656), (50600,-0.404161), (50601,-0.145847), (50602,0.097139), (50603,0.023340), (50604,-0.139637), (50605,-0.107068), (50606,-0.293739), (50607,-0.333161), (50608,-0.493358), (50609,-0.208563), (50610,0.005162), (50611,0.008470), (50612,-0.140112), (50613,-0.023468), (50614,-0.042921), (50615,-0.098135), (50616,-0.509156), (50617,-0.215544), (50618,0.025125), (50619,0.006598), (50620,-0.142447), (50621,-0.162827), (50622,-0.399197), (50623,-0.443265), (50624,-0.597889), (50625,-0.327496), (50626,-0.056639), (50627,-0.130438), (50628,-0.344510), (50629,-0.152156), (50630,-0.196687), (50631,-0.241225), (50632,-0.349394), (50633,-0.069708), (50634,0.159809), (50635,0.137569), (50636,-0.028201), (50637,-0.034649), (50638,-0.218064), (50639,-0.245877), (50640,-0.421866), (50641,-0.154722), (50642,0.093836), (50643,0.039549), (50644,-0.124361), (50645,0.032696), (50646,-0.011841), (50647,-0.084243), (50648,-0.500837), (50649,-0.175635), (50650,-0.005573), (50651,-0.035709), (50652,-0.152243), (50653,-0.178196), (50654,-0.346752), (50655,-0.402430), (50656,-0.564950), (50657,-0.298270), (50658,-0.075258), (50659,-0.117936), (50660,-0.260475), (50661,-0.101565), (50662,-0.172107), (50663,-0.204103), (50664,-0.355471), (50665,-0.091584), (50666,0.154658), (50667,0.070178), (50668,-0.046820), (50669,-0.032367), (50670,-0.221355), (50671,-0.290977), (50672,-0.465569), (50673,-0.201212), (50674,0.036664), (50675,-0.023665), (50676,-0.158772), (50677,-0.004508), (50678,-0.067154), (50679,-0.131660), (50680,-0.186880), (50681,0.082580), (50682,-0.027912), (50683,0.303333), (50684,0.149641), (50685,0.172461), (50686,0.024806), (50687,-0.079650), (50688,-0.185959), (50689,0.062600), (50690,-0.072049), (50691,0.262908), (50692,0.073456), (50693,0.253732), (50694,0.111656), (50695,0.098239), (50696,-0.191080), (50697,0.109037), (50698,-0.042331), (50699,0.304242), (50700,0.145905), (50701,0.164541), (50702,-0.003082), (50703,-0.050870), (50704,-0.234291), (50705,0.037035), (50706,-0.112016), (50707,0.231307), (50708,0.031167), (50709,0.213765), (50710,0.089804), (50711,0.114947), (50712,0.171666), (50713,-0.029864), (50714,-0.121777), (50715,0.129105), (50716,0.186294), (50717,0.032603), (50718,-0.021221), (50719,-0.207892), (50720,0.088975), (50721,-0.107445), (50722,-0.167775), (50723,0.084040), (50724,0.217409), (50725,0.093442), (50726,0.045191), (50727,-0.068550), (50728,-0.017867), (50729,-0.147400), (50730,0.194990), (50731,0.065913), (50732,0.100805), (50733,-0.067745), (50734,-0.177310), (50735,-0.293375), (50736,-0.018805), (50737,-0.170636), (50738,0.154565), (50739,0.047323), (50740,0.176046), (50741,0.010739), (50742,0.035418), (50743,-0.134065), (50744,0.171626), (50745,0.005399), (50746,-0.038676), (50747,0.186195), (50748,0.187650), (50749,0.028849), (50750,0.025651), (50751,-0.147082), (50752,0.158145), (50753,-0.046172), (50754,-0.139482), (50755,0.117443), (50756,0.248489), (50757,0.111516), (50758,0.036791), (50759,-0.036080), (50760,0.146061), (50761,0.040215), (50762,-0.022901), (50763,0.205220), (50764,0.230362), (50765,0.106395), (50766,0.017274), (50767,-0.150819), (50768,0.133507), (50769,-0.043409), (50770,-0.092586), (50771,0.142504), (50772,0.327895), (50773,0.167704), (50774,0.087400), (50775,0.009888), (50776,0.203175), (50777,0.017430), (50778,0.008666), (50779,0.252115), (50780,0.246137), (50781,0.103128), (50782,0.050694), (50783,-0.128544), (50784,0.137666), (50785,0.000700), (50786,-0.077745), (50787,0.193582), (50788,0.337163), (50789,0.148169), (50790,0.088309), (50791,0.014511), (50792,0.120009), (50793,-0.060156), (50794,0.273868), (50795,0.139225), (50796,0.145319), (50797,-0.019054), (50798,-0.110505), (50799,-0.242831), (50800,0.033135), (50801,-0.116373), (50802,0.246455), (50803,0.056997), (50804,0.183860), (50805,0.046894), (50806,0.067384), (50807,-0.070045), (50808,-0.007746), (50809,-0.172590), (50810,0.165624), (50811,-0.003396), (50812,0.023600), (50813,-0.112903), (50814,-0.234547), (50815,-0.398920), (50816,-0.253479), (50817,-0.430858), (50818,-0.048982), (50819,-0.191064), (50820,-0.029361), (50821,-0.201630), (50822,-0.145837), (50823,-0.291632), (50824,-0.437890), (50825,-0.159138), (50826,0.088957), (50827,0.037920), (50828,-0.130630), (50829,-0.138474), (50830,-0.294952), (50831,-0.335306), (50832,-0.498747), (50833,-0.204202), (50834,-0.005343), (50835,-0.013644), (50836,-0.215644), (50837,-0.074848), (50838,-0.185804), (50839,-0.203861), (50840,-0.343156), (50841,-0.051861), (50842,-0.193937), (50843,0.121979), (50844,-0.003379), (50845,-0.022369), (50846,-0.167700), (50847,-0.206659), (50848,-0.374752), (50849,-0.067659), (50850,-0.231569), (50851,0.074121), (50852,-0.077710), (50853,0.056586), (50854,-0.123116), (50855,-0.067787), (50856,-0.380800), (50857,-0.112266), (50858,0.138159), (50859,0.077366), (50860,-0.075399), (50861,-0.077664), (50862,-0.249933), (50863,-0.294008), (50864,-0.450949), (50865,-0.156867), (50866,0.047102), (50867,0.012326), (50868,-0.116280), (50869,0.049136), (50870,-0.020486), (50871,-0.072450), (50872,-0.490903), (50873,-0.244198), (50874,-0.022114), (50875,-0.058286), (50876,-0.166461), (50877,-0.135746), (50878,-0.362830), (50879,-0.399002), (50880,-0.581490), (50881,-0.280440), (50882,0.010855), (50883,-0.076876), (50884,-0.302100), (50885,-0.114386), (50886,-0.211409), (50887,-0.248514), (50888,-0.454691), (50889,-0.144354), (50890,0.079590), (50891,0.037375), (50892,-0.125138), (50893,-0.131586), (50894,-0.305252), (50895,-0.363722), (50896,-0.515553), (50897,-0.244697), (50898,0.010368), (50899,-0.033700), (50900,-0.172989), (50901,-0.060528), (50902,-0.117602), (50903,-0.150060), (50904,-0.337658), (50905,-0.039864), (50906,-0.167075), (50907,0.135829), (50908,-0.038763), (50909,-0.000152), (50910,-0.171032), (50911,-0.270841), (50912,-0.395271), (50913,-0.115586), (50914,-0.245126), (50915,0.072186), (50916,-0.082438), (50917,0.083911), (50918,-0.082322), (50919,-0.059509), (50920,-0.223882), (50921,0.033969), (50922,-0.124832), (50923,0.216168), (50924,0.057367), (50925,0.069968), (50926,-0.080937), (50927,-0.158918), (50928,-0.325152), (50929,-0.045003), (50930,-0.181505), (50931,0.158092), (50932,0.028558), (50933,0.176786), (50934,0.043996), (50935,0.080285), (50936,-0.082229), (50937,0.157970), (50938,0.002419), (50939,0.338773), (50940,0.161857), (50941,0.203718), (50942,-0.004318), (50943,-0.059538), (50944,-0.237380), (50945,0.046945), (50946,-0.131360), (50947,0.223102), (50948,0.072197), (50949,0.212536), (50950,0.021681), (50951,0.076084), (50952,-0.218814), (50953,0.057152), (50954,-0.105825), (50955,0.250497), (50956,0.119104), (50957,0.112193), (50958,-0.047071), (50959,-0.106004), (50960,-0.283853), (50961,0.006515), (50962,-0.162041), (50963,0.132973), (50964,0.001110), (50965,0.177215), (50966,0.042566), (50967,0.065848), (50968,0.122105), (50969,-0.003716), (50970,-0.070545), (50971,0.148290), (50972,0.185041), (50973,0.032277), (50974,-0.025723), (50975,-0.204499), (50976,0.053352), (50977,-0.100339), (50978,-0.162058), (50979,0.106938), (50980,0.220796), (50981,0.092653), (50982,0.039292), (50983,-0.041006), (50984,0.144385), (50985,-0.048792), (50986,-0.114225), (50987,0.130151), (50988,0.100948), (50989,-0.006757), (50990,-0.073123), (50991,-0.229600), (50992,0.055189), (50993,-0.118477), (50994,-0.147217), (50995,0.082300), (50996,0.223565), (50997,0.033644), (50998,0.003045), (50999,-0.057748), (51000,0.143898), (51001,-0.013042), (51002,-0.087774), (51003,0.163578), (51004,0.147844), (51005,0.044315), (51006,-0.021588), (51007,-0.182711), (51008,0.115089), (51009,-0.023273), (51010,-0.084993), (51011,0.121763), (51012,0.271387), (51013,0.059632), (51014,0.026709), (51015,-0.068454), (51016,0.133192), (51017,-0.021425), (51018,-0.079432), (51019,0.163091), (51020,0.195202), (51021,0.101429), (51022,0.022058), (51023,-0.154858), (51024,0.134114), (51025,-0.051161), (51026,-0.124033), (51027,0.117563), (51028,0.282052), (51029,0.099094), (51030,0.010900), (51031,-0.059185), (51032,0.155473), (51033,0.008745), (51034,-0.033000), (51035,0.187225), (51036,0.244414), (51037,0.074931), (51038,0.040619), (51039,-0.122828), (51040,0.120621), (51041,-0.038643), (51042,-0.084570), (51043,0.150056), (51044,0.288535), (51045,0.122765), (51046,0.062435), (51047,0.005825), (51048,0.093209), (51049,-0.071165), (51050,0.286554), (51051,0.122643), (51052,0.138493), (51053,0.006630), (51054,-0.089929), (51055,-0.225969), (51056,0.090410), (51057,-0.053988), (51058,0.298621), (51059,0.111949), (51060,0.236026), (51061,0.054927), (51062,0.126519), (51063,-0.014630), (51064,-0.056381), (51065,-0.197067), (51066,0.122562), (51067,-0.003259), (51068,0.009805), (51069,-0.160605), (51070,-0.236726), (51071,-0.406673), (51072,-0.065216), (51073,-0.262106), (51074,-0.352623), (51075,-0.059005), (51076,0.067394), (51077,-0.087693), (51078,-0.118292), (51079,-0.179085), (51080,-0.484202), (51081,-0.191511), (51082,0.059834), (51083,0.029704), (51084,-0.143498), (51085,-0.111393), (51086,-0.262297), (51087,-0.340736), (51088,-0.490250), (51089,-0.189200), (51090,0.038457), (51091,-0.009324), (51092,-0.172307), (51093,-0.025933), (51094,-0.139217), (51095,-0.221838), (51096,-0.336043), (51097,-0.047072), (51098,-0.192867), (51099,0.187606), (51100,0.017660), (51101,0.041406), (51102,-0.120644), (51103,-0.188870), (51104,-0.347671), (51105,-0.087033), (51106,-0.259302), (51107,0.074728), (51108,-0.062708), (51109,0.106428), (51110,-0.059805), (51111,-0.018408), (51112,-0.439647), (51113,-0.198521), (51114,0.072335), (51115,-0.013999), (51116,-0.170013), (51117,-0.164846), (51118,-0.345481), (51119,-0.391408), (51120,-0.559032), (51121,-0.271920), (51122,0.017052), (51123,-0.023303), (51124,-0.213224), (51125,-0.034802), (51126,-0.128569), (51127,-0.156382), (51128,-0.371387), (51129,-0.053155), (51130,-0.215669), (51131,0.071443), (51132,-0.052054), (51133,-0.065465), (51134,-0.162951), (51135,-0.212599), (51136,-0.403446), (51137,-0.119121), (51138,-0.251447), (51139,0.025915), (51140,-0.136135), (51141,0.039500), (51142,-0.122087), (51143,-0.085799), (51144,-0.433652), (51145,-0.099621), (51146,0.115957), (51147,0.048665), (51148,-0.123142), (51149,-0.083604), (51150,-0.254013), (51151,-0.328745), (51152,-0.508447), (51153,-0.237590), (51154,0.050918), (51155,0.006850), (51156,-0.169139), (51157,0.021362), (51158,-0.055223), (51159,-0.113693), (51160,-0.315687), (51161,-0.049940), (51162,-0.198521), (51163,0.132253), (51164,-0.016792), (51165,-0.006051), (51166,-0.129549), (51167,-0.192201), (51168,-0.356111), (51169,-0.065280), (51170,-0.265420), (51171,0.095548), (51172,-0.090660), (51173,0.069183), (51174,-0.084971), (51175,-0.051933), (51176,-0.199124), (51177,0.065696), (51178,-0.057338), (51179,0.259041), (51180,0.106740), (51181,0.135132), (51182,-0.015773), (51183,-0.110936), (51184,-0.257658), (51185,0.000657), (51186,-0.136779), (51187,0.173564), (51188,0.039378), (51189,0.178320), (51190,0.051573), (51191,0.070209), (51192,-0.146656), (51193,0.099586), (51194,-0.054569), (51195,0.345416), (51196,0.182433), (51197,0.186674), (51198,0.018117), (51199,-0.066827), (51200,-0.503395), (51201,-0.653837), (51202,0.020203), (51203,-0.122343), (51204,-0.196141), (51205,-0.293158), (51206,-0.046922), (51207,-0.232660), (51208,-0.457421), (51209,-0.576273), (51210,0.050848), (51211,-0.076362), (51212,-0.142734), (51213,-0.272731), (51214,-0.242949), (51215,-0.436120), (51216,-0.477408), (51217,-0.633416), (51218,0.048050), (51219,-0.094952), (51220,-0.185939), (51221,-0.306187), (51222,-0.074810), (51223,-0.202953), (51224,-0.391484), (51225,-0.107622), (51226,-0.238552), (51227,0.117306), (51228,-0.041958), (51229,-0.076270), (51230,-0.237394), (51231,-0.315375), (51232,-0.441658), (51233,-0.151760), (51234,-0.333316), (51235,0.015574), (51236,-0.127435), (51237,-0.023333), (51238,-0.152866), (51239,-0.127261), (51240,-0.501588), (51241,-0.198215), (51242,0.048484), (51243,-0.009516), (51244,-0.223595), (51245,-0.194276), (51246,-0.412994), (51247,-0.454276), (51248,-0.594961), (51249,-0.344080), (51250,-0.073223), (51251,-0.119151), (51252,-0.283988), (51253,-0.131577), (51254,-0.219777), (51255,-0.245730), (51256,-0.561993), (51257,-0.278594), (51258,-0.054187), (51259,-0.139601), (51260,-0.277030), (51261,-0.273259), (51262,-0.436706), (51263,-0.468232), (51264,-0.661403), (51265,-0.393332), (51266,-0.128518), (51267,-0.203707), (51268,-0.357861), (51269,-0.185482), (51270,-0.262530), (51271,-0.314494), (51272,-0.511848), (51273,-0.264679), (51274,-0.083008), (51275,-0.150300), (51276,-0.252433), (51277,-0.229150), (51278,-0.393060), (51279,-0.441311), (51280,-0.614977), (51281,-0.332968), (51282,-0.118780), (51283,-0.116868), (51284,-0.265450), (51285,-0.126045), (51286,-0.218885), (51287,-0.282464), (51288,-0.366945), (51289,-0.112814), (51290,-0.323636), (51291,0.078672), (51292,-0.060617), (51293,-0.033158), (51294,-0.181270), (51295,-0.244850), (51296,-0.405973), (51297,-0.138830), (51298,-0.295777), (51299,0.037790), (51300,-0.092676), (51301,0.057875), (51302,-0.093957), (51303,-0.066961), (51304,-0.354427), (51305,-0.497435), (51306,0.148270), (51307,-0.011457), (51308,-0.068067), (51309,-0.200857), (51310,-0.204055), (51311,-0.372605), (51312,-0.454769), (51313,-0.564798), (51314,0.110638), (51315,-0.044913), (51316,-0.107559), (51317,-0.261250), (51318,-0.010831), (51319,-0.166382), (51320,-0.477072), (51321,-0.202496), (51322,0.013546), (51323,-0.019377), (51324,-0.162849), (51325,-0.147925), (51326,-0.331347), (51327,-0.398640), (51328,-0.789686), (51329,-0.539730), (51330,-0.256801), (51331,-0.374726), (51332,-0.429940), (51333,-0.523713), (51334,-0.360620), (51335,-0.500835), (51336,-0.639668), (51337,-0.393426), (51338,-0.145330), (51339,-0.294839), (51340,-0.358881), (51341,-0.523255), (51342,-0.476754), (51343,-0.647164), (51344,-0.725145), (51345,-0.481689), (51346,-0.155561), (51347,-0.350592), (51348,-0.398373), (51349,-0.489823), (51350,-0.354137), (51351,-0.495286), (51352,-0.664769), (51353,-0.443612), (51354,-0.134665), (51355,-0.266991), (51356,-0.325925), (51357,-0.465214), (51358,-0.536226), (51359,-0.686667), (51360,-0.701474), (51361,-0.443623), (51362,-0.180199), (51363,-0.359901), (51364,-0.397470), (51365,-0.441074), (51366,-0.302132), (51367,-0.447928), (51368,-0.529159), (51369,-0.266198), (51370,0.007915), (51371,-0.129521), (51372,-0.185668), (51373,-0.407173), (51374,-0.418730), (51375,-0.594250), (51376,-0.642037), (51377,-0.376753), (51378,-0.089178), (51379,-0.289782), (51380,-0.306912), (51381,-0.367242), (51382,-0.197179), (51383,-0.353657), (51384,-0.691284), (51385,-0.478956), (51386,-0.162113), (51387,-0.337169), (51388,-0.357549), (51389,-0.536788), (51390,-0.514438), (51391,-0.709932), (51392,-0.777688), (51393,-0.543531), (51394,-0.233189), (51395,-0.454700), (51396,-0.505737), (51397,-0.543769), (51398,-0.401577), (51399,-0.556658), (51400,-0.611415), (51401,-0.359137), (51402,-0.048794), (51403,-0.199236), (51404,-0.223335), (51405,-0.450413), (51406,-0.441996), (51407,-0.613338), (51408,-0.696893), (51409,-0.385623), (51410,-0.109187), (51411,-0.303755), (51412,-0.363621), (51413,-0.476899), (51414,-0.315196), (51415,-0.452168), (51416,-0.739634), (51417,-0.435797), (51418,-0.168654), (51419,-0.360435), (51420,-0.356200), (51421,-0.527543), (51422,-0.532131), (51423,-0.752240), (51424,-0.767980), (51425,-0.512452), (51426,-0.242985), (51427,-0.407822), (51428,-0.479297), (51429,-0.508970), (51430,-0.342157), (51431,-0.514896), (51432,-0.565470), (51433,-0.256061), (51434,-0.420434), (51435,-0.098482), (51436,-0.280507), (51437,-0.380317), (51438,-0.485236), (51439,-0.449874), (51440,-0.631899), (51441,-0.314130), (51442,-0.475254), (51443,-0.203001), (51444,-0.347400), (51445,-0.313441), (51446,-0.457840), (51447,-0.342586), (51448,-0.377368), (51449,-0.506438), (51450,0.157846), (51451,0.006008), (51452,-0.025981), (51453,-0.197324), (51454,-0.215381), (51455,-0.386260), (51456,-0.451700), (51457,-0.570087), (51458,0.091410), (51459,-0.036270), (51460,-0.065943), (51461,-0.256327), (51462,-0.038419), (51463,-0.152630), (51464,-0.362063), (51465,-0.431679), (51466,-0.145957), (51467,0.125363), (51468,-0.075704), (51469,-0.113735), (51470,-0.281359), (51471,-0.266442), (51472,-0.410377), (51473,-0.501827), (51474,-0.253262), (51475,0.054751), (51476,-0.127274), (51477,-0.156477), (51478,-0.203338), (51479,-0.071365), (51480,-0.446156), (51481,-0.190158), (51482,0.043999), (51483,0.031051), (51484,-0.169089), (51485,-0.156952), (51486,-0.342233), (51487,-0.409062), (51488,-0.562290), (51489,-0.257520), (51490,-0.028936), (51491,-0.064645), (51492,-0.193252), (51493,-0.079858), (51494,-0.139254), (51495,-0.186578), (51496,-0.505627), (51497,-0.262642), (51498,0.036549), (51499,-0.195638), (51500,-0.214165), (51501,-0.401763), (51502,-0.383590), (51503,-0.531245), (51504,-0.582282), (51505,-0.332790), (51506,-0.079585), (51507,-0.218411), (51508,-0.272698), (51509,-0.321419), (51510,-0.183404), (51511,-0.369148), (51512,-0.476384), (51513,-0.149323), (51514,0.107132), (51515,0.046339), (51516,-0.103632), (51517,-0.113800), (51518,-0.276777), (51519,-0.357081), (51520,-0.527954), (51521,-0.229690), (51522,0.002613), (51523,-0.029382), (51524,-0.221163), (51525,-0.038095), (51526,-0.123040), (51527,-0.123915), (51528,-0.329628), (51529,-0.499574), (51530,0.164710), (51531,0.008696), (51532,-0.015867), (51533,-0.165839), (51534,-0.149062), (51535,-0.305077), (51536,-0.405813), (51537,-0.556717), (51538,0.161912), (51539,0.021226), (51540,-0.036781), (51541,-0.177930), (51542,0.104542), (51543,-0.129968), (51544,-0.371454), (51545,-0.107560), (51546,0.124743), (51547,0.069986), (51548,-0.111106), (51549,-0.069708), (51550,-0.260562), (51551,-0.296734), (51552,-0.457395), (51553,-0.176783), (51554,0.078282), (51555,0.010990), (51556,-0.154780), (51557,0.009246), (51558,-0.096606), (51559,-0.129065), (51560,-0.382154), (51561,-0.150777), (51562,0.144231), (51563,-0.043367), (51564,-0.106947), (51565,-0.270393), (51566,-0.265689), (51567,-0.428209), (51568,-0.452766), (51569,-0.236254), (51570,0.064790), (51571,-0.070317), (51572,-0.132506), (51573,-0.186793), (51574,-0.048314), (51575,-0.226163), (51576,-0.578656), (51577,-0.328701), (51578,-0.017431), (51579,-0.203176), (51580,-0.250964), (51581,-0.459926), (51582,-0.428285), (51583,-0.604737), (51584,-0.898702), (51585,-0.191219), (51586,-0.341197), (51587,-0.410349), (51588,-0.515268), (51589,-0.287147), (51590,-0.497507), (51591,-0.509521), (51592,-0.640457), (51593,-0.448097), (51594,-0.139614), (51595,-0.269617), (51596,-0.324374), (51597,-0.475272), (51598,-0.512841), (51599,-0.634948), (51600,-0.685985), (51601,-0.469937), (51602,-0.162387), (51603,-0.300749), (51604,-0.371298), (51605,-0.440914), (51606,-0.293149), (51607,-0.488643), (51608,-0.498341), (51609,-0.639490), (51610,0.062420), (51611,-0.107532), (51612,-0.208268), (51613,-0.336875), (51614,-0.338214), (51615,-0.520239), (51616,-0.599147), (51617,-0.765380), (51618,-0.054641), (51619,-0.211588), (51620,-0.212920), (51621,-0.400988), (51622,-0.180293), (51623,-0.331661), (51624,-0.549917), (51625,-0.303681), (51626,-0.024928), (51627,-0.178620), (51628,-0.213395), (51629,-0.387524), (51630,-0.380967), (51631,-0.569961), (51632,-0.615889), (51633,-0.395194), (51634,-0.124338), (51635,-0.256664), (51636,-0.290976), (51637,-0.311357), (51638,-0.199822), (51639,-0.340044), (51640,-0.689751), (51641,-0.463020), (51642,-0.161043), (51643,-0.352361), (51644,-0.405721), (51645,-0.580777), (51646,-0.554708), (51647,-0.705612), (51648,-0.758509), (51649,-0.516450), (51650,-0.242807), (51651,-0.358872), (51652,-0.434530), (51653,-0.543162), (51654,-0.412116), (51655,-0.553265), (51656,-0.623814), (51657,-0.396157), (51658,-0.093710), (51659,-0.234859), (51660,-0.303548), (51661,-0.506474), (51662,-0.455791), (51663,-0.607622), (51664,-0.674921), (51665,-0.439361), (51666,-0.131811), (51667,-0.306404), (51668,-0.326321), (51669,-0.434489), (51670,-0.287651), (51671,-0.445989), (51672,-0.533719), (51673,-0.666972), (51674,0.024249), (51675,-0.159172), (51676,-0.227855), (51677,-0.360181), (51678,-0.364769), (51679,-0.500809), (51680,-0.576930), (51681,-0.730158), (51682,-0.079343), (51683,-0.241394), (51684,-0.307759), (51685,-0.453091), (51686,-0.199423), (51687,-0.309915), (51688,-0.403218), (51689,-0.554123), (51690,0.142678), (51691,-0.025879), (51692,-0.104787), (51693,-0.250118), (51694,-0.239378), (51695,-0.406075), (51696,-0.480800), (51697,-0.628454), (51698,-0.010620), (51699,-0.159665), (51700,-0.202806), (51701,-0.354637), (51702,-0.101896), (51703,-0.255587), (51704,-0.347500), (51705,-0.502118), (51706,0.165879), (51707,0.013121), (51708,-0.017485), (51709,-0.189291), (51710,-0.215707), (51711,-0.380081), (51712,-0.396284), (51713,-0.575053), (51714,0.082261), (51715,-0.057498), (51716,-0.139192), (51717,-0.250147), (51718,-0.028526), (51719,-0.196150), (51720,-0.402332), (51721,-0.588534), (51722,0.077140), (51723,-0.048217), (51724,-0.115973), (51725,-0.276170), (51726,-0.269612), (51727,-0.411688), (51728,-0.491986), (51729,-0.636855), (51730,0.055763), (51731,-0.054265), (51732,-0.135496), (51733,-0.250634), (51734,-0.037836), (51735,-0.196173), (51736,-0.452518), (51737,-0.190021), (51738,0.078513), (51739,0.024226), (51740,-0.129002), (51741,-0.174466), (51742,-0.362065), (51743,-0.352720), (51744,-0.529636), (51745,-0.275962), (51746,-0.053877), (51747,-0.066825), (51748,-0.249783), (51749,-0.104335), (51750,-0.175347), (51751,-0.227317), (51752,-0.525465), (51753,-0.227201), (51754,0.014858), (51755,0.020489), (51756,-0.154104), (51757,-0.167521), (51758,-0.375087), (51759,-0.455392), (51760,-0.614656), (51761,-0.342872), (51762,-0.051578), (51763,-0.102145), (51764,-0.257233), (51765,-0.128973), (51766,-0.179547), (51767,-0.225011), (51768,-0.500868), (51769,-0.190062), (51770,-0.006530), (51771,-0.055244), (51772,-0.209862), (51773,-0.205164), (51774,-0.349563), (51775,-0.385272), (51776,-0.512489), (51777,-0.273216), (51778,-0.058101), (51779,-0.109138), (51780,-0.230312), (51781,-0.079761), (51782,-0.157273), (51783,-0.196231), (51784,-0.471154), (51785,-0.172897), (51786,0.083101), (51787,0.004656), (51788,-0.181088), (51789,-0.136904), (51790,-0.315673), (51791,-0.368570), (51792,-0.534340), (51793,-0.228644), (51794,0.014342), (51795,-0.058060), (51796,-0.243341), (51797,-0.069559), (51798,-0.122920), (51799,-0.188822), (51800,-0.452600), (51801,-0.166414), (51802,0.058463), (51803,0.016711), (51804,-0.147662), (51805,-0.140171), (51806,-0.327776), (51807,-0.392745), (51808,-0.530181), (51809,-0.234240), (51810,-0.000540), (51811,-0.041358), (51812,-0.185294), (51813,-0.040316), (51814,-0.101109), (51815,-0.171194), (51816,-0.506962), (51817,0.186119), (51818,-0.011234), (51819,-0.082246), (51820,-0.271241), (51821,-0.255391), (51822,-0.369133), (51823,-0.455936), (51824,-0.605914), (51825,0.091813), (51826,-0.077200), (51827,-0.126384), (51828,-0.294471), (51829,-0.030120), (51830,-0.227011), (51831,-0.270152), (51832,-0.706251), (51833,-0.006670), (51834,-0.145959), (51835,-0.202106), (51836,-0.367876), (51837,-0.332051), (51838,-0.456481), (51839,-0.521451), (51840,-0.650991), (51841,-0.406608), (51842,-0.173372), (51843,-0.295479), (51844,-0.349303), (51845,-0.446326), (51846,-0.290665), (51847,-0.443423), (51848,-0.612443), (51849,-0.335087), (51850,-0.091168), (51851,-0.263437), (51852,-0.283354), (51853,-0.434722), (51854,-0.462071), (51855,-0.603220), (51856,-0.652404), (51857,-0.400589), (51858,-0.141812), (51859,-0.285747), (51860,-0.360009), (51861,-0.433344), (51862,-0.269781), (51863,-0.435088), (51864,-0.653806), (51865,-0.307233), (51866,-0.445133), (51867,-0.157088), (51868,-0.328430), (51869,-0.407802), (51870,-0.555457), (51871,-0.544253), (51872,-0.655671), (51873,-0.318861), (51874,-0.499026), (51875,-0.196116), (51876,-0.387433), (51877,-0.355328), (51878,-0.491831), (51879,-0.367291), (51880,-0.338435), (51881,-0.389473), (51882,-0.509257), (51883,-0.239327), (51884,-0.426925), (51885,-0.517442), (51886,-0.652555), (51887,-0.654820), (51888,-0.404865), (51889,-0.410849), (51890,-0.563607), (51891,-0.289501), (51892,-0.361440), (51893,-0.418519), (51894,-0.611690), (51895,-0.467176), (51896,-0.625513), (51897,-0.278940), (51898,-0.434491), (51899,-0.162238), (51900,-0.295491), (51901,-0.355820), (51902,-0.511835), (51903,-0.523855), (51904,-0.668254), (51905,-0.347699), (51906,-0.483275), (51907,-0.191980), (51908,-0.341488), (51909,-0.329358), (51910,-0.486299), (51911,-0.350143), (51912,-0.525663), (51913,-0.206034), (51914,-0.377840), (51915,-0.114879), (51916,-0.234200), (51917,-0.369313), (51918,-0.490024), (51919,-0.479283), (51920,-0.635297), (51921,-0.277579), (51922,-0.414082), (51923,-0.162273), (51924,-0.292270), (51925,-0.289426), (51926,-0.449623), (51927,-0.282810), (51928,-0.675252), (51929,-0.312424), (51930,-0.448934), (51931,-0.180863), (51932,-0.339194), (51933,-0.424608), (51934,-0.561111), (51935,-0.555480), (51936,-0.674801), (51937,-0.352849), (51938,-0.499108), (51939,-0.225465), (51940,-0.354998), (51941,-0.305241), (51942,-0.457072), (51943,-0.313491), (51944,-0.496443), (51945,-0.161022), (51946,-0.324469), (51947,-0.072191), (51948,-0.221699), (51949,-0.327081), (51950,-0.490065), (51951,-0.474215), (51952,-0.613040), (51953,-0.272510), (51954,-0.422018), (51955,-0.151162), (51956,-0.305786), (51957,-0.265779), (51958,-0.431085), (51959,-0.291216), (51960,-0.483924), (51961,-0.132705), (51962,-0.324486), (51963,-0.050380), (51964,-0.179450), (51965,-0.242566), (51966,-0.420871), (51967,-0.413387), (51968,-0.552213), (51969,-0.234907), (51970,-0.360728), (51971,-0.038313), (51972,-0.201759), (51973,-0.147820), (51974,-0.315443), (51975,-0.202518), (51976,-0.520635), (51977,-0.186147), (51978,-0.342155), (51979,-0.081517), (51980,-0.215703), (51981,-0.288569), (51982,-0.467344), (51983,-0.482151), (51984,-0.626087), (51985,-0.274874), (51986,-0.400231), (51987,-0.156312), (51988,-0.317899), (51989,-0.281611), (51990,-0.451094), (51991,-0.294507), (51992,-0.410572), (51993,-0.560080), (51994,0.109313), (51995,-0.033695), (51996,-0.093098), (51997,-0.236101), (51998,-0.249054), (51999,-0.400886), (52000,-0.464928), (52001,-0.612583), (52002,0.055883), (52003,-0.112210), (52004,-0.174393), (52005,-0.340163), (52006,-0.094384), (52007,-0.246215), (52008,-0.587099), (52009,-0.310670), (52010,-0.024485), (52011,-0.200474), (52012,-0.247328), (52013,-0.421457), (52014,-0.392602), (52015,-0.546756), (52016,-0.611732), (52017,-0.392428), (52018,-0.060726), (52019,-0.234386), (52020,-0.282637), (52021,-0.388025), (52022,-0.251406), (52023,-0.400451), (52024,-0.515589), (52025,-0.318120), (52026,-0.051446), (52027,-0.177730), (52028,-0.219011), (52029,-0.410329), (52030,-0.358249), (52031,-0.551420), (52032,-0.590848), (52033,-0.330210), (52034,-0.064926), (52035,-0.190747), (52036,-0.253400), (52037,-0.323942), (52038,-0.187323), (52039,-0.329405), (52040,-0.492382), (52041,-0.206197), (52042,0.092061), (52043,-0.106683), (52044,-0.166080), (52045,-0.361110), (52046,-0.335041), (52047,-0.483623), (52048,-0.558818), (52049,-0.329301), (52050,-0.034287), (52051,-0.177295), (52052,-0.273855), (52053,-0.323032), (52054,-0.155293), (52055,-0.339641), (52056,-0.368850), (52057,-0.497457), (52058,0.132456), (52059,0.010812), (52060,-0.043938), (52061,-0.197166), (52062,-0.223119), (52063,-0.390748), (52064,-0.469193), (52065,-0.652608), (52066,0.068344), (52067,-0.088134), (52068,-0.129885), (52069,-0.308654), (52070,-0.051266), (52071,-0.179410), (52072,-0.175175), (52073,-0.361383), (52074,-0.055687), (52075,-0.208914), (52076,-0.269238), (52077,-0.414569), (52078,-0.417768), (52079,-0.529186), (52080,-0.204911), (52081,-0.365571), (52082,-0.058022), (52083,-0.260015), (52084,-0.227447), (52085,-0.330969), (52086,-0.228263), (52087,-0.373126), (52088,-0.531926), (52089,-0.223913), (52090,0.048340), (52091,-0.118820), (52092,-0.189832), (52093,-0.366748), (52094,-0.359727), (52095,-0.508302), (52096,-0.655493), (52097,-0.702817), (52098,-0.473764), (52099,-0.214053), (52100,-0.370530), (52101,-0.391844), (52102,-0.466569), (52103,-0.295110), (52104,-0.704277), (52105,-0.350272), (52106,-0.520225), (52107,-0.258191), (52108,-0.376115), (52109,-0.442481), (52110,-0.625433), (52111,-0.607729), (52112,-0.769780), (52113,-0.382801), (52114,-0.550424), (52115,-0.274921), (52116,-0.457410), (52117,-0.413226), (52118,-0.562740), (52119,-0.362021), (52120,-0.546832), (52121,-0.587187), (52122,-0.380431), (52123,-0.080771), (52124,-0.247467), (52125,-0.319412), (52126,-0.473104), (52127,-0.468399), (52128,-0.623950), (52129,-0.679164), (52130,-0.412490), (52131,-0.146743), (52132,-0.324585), (52133,-0.374696), (52134,-0.438275), (52135,-0.260780), (52136,-0.631388), (52137,-0.329875), (52138,-0.406923), (52139,-0.590808), (52140,-0.261423), (52141,-0.461563), (52142,-0.499132), (52143,-0.656073), (52144,-0.673666), (52145,-0.421858), (52146,-0.432019), (52147,-0.613581), (52148,-0.354333), (52149,-0.393298), (52150,-0.442012), (52151,-0.613818), (52152,-0.567774), (52153,-0.642036), (52154,-0.421348), (52155,-0.117042), (52156,-0.272593), (52157,-0.350104), (52158,-0.531666), (52159,-0.487945), (52160,-0.670903), (52161,-0.711258), (52162,-0.497997), (52163,-0.194623), (52164,-0.357143), (52165,-0.397028), (52166,-0.472223), (52167,-0.320739), (52168,-0.546427), (52169,-0.322952), (52170,-0.388385), (52171,-0.560191), (52172,-0.283298), (52173,-0.455105), (52174,-0.498246), (52175,-0.650541), (52176,-0.638410), (52177,-0.400527), (52178,-0.407439), (52179,-0.571812), (52180,-0.327436), (52181,-0.418417), (52182,-0.429047), (52183,-0.602707), (52184,-0.603119), (52185,-0.621639), (52186,-0.392585), (52187,-0.128235), (52188,-0.237330), (52189,-0.299519), (52190,-0.502909), (52191,-0.502851), (52192,-0.680700), (52193,-0.711299), (52194,-0.466917), (52195,-0.169586), (52196,-0.307948), (52197,-0.327395), (52198,-0.417455), (52199,-0.271544), (52200,-0.361135), (52201,-0.512503), (52202,-0.126913), (52203,-0.287574), (52204,-0.009285), (52205,-0.167622), (52206,-0.245133), (52207,-0.459675), (52208,-0.441966), (52209,-0.582188), (52210,-0.235615), (52211,-0.366082), (52212,-0.093372), (52213,-0.229411), (52214,-0.238176), (52215,-0.332412), (52216,-0.375090), (52217,-0.428914), (52218,-0.169203), (52219,0.107690), (52220,-0.072476), (52221,-0.136988), (52222,-0.317617), (52223,-0.320345), (52224,-0.432234), (52225,-0.473052), (52226,-0.231926), (52227,0.058442), (52228,-0.110577), (52229,-0.160682), (52230,-0.234950), (52231,-0.049559), (52232,-0.284533), (52233,-0.446583), (52234,-0.102340), (52235,-0.275536), (52236,-0.022331), (52237,-0.161626), (52238,-0.247961), (52239,-0.392829), (52240,-0.418319), (52241,-0.552035), (52242,-0.210115), (52243,-0.376342), (52244,-0.118027), (52245,-0.294016), (52246,-0.234040), (52247,-0.399804), (52248,-0.589262), (52249,-0.662133), (52250,-0.420074), (52251,-0.125993), (52252,-0.272715), (52253,-0.272193), (52254,-0.434707), (52255,-0.433722), (52256,-0.599029), (52257,-0.650993), (52258,-0.397788), (52259,-0.103707), (52260,-0.235100), (52261,-0.342806), (52262,-0.403135), (52263,-0.233999), (52264,-0.409525), (52265,-0.469848), (52266,-0.241728), (52267,0.047707), (52268,-0.111093), (52269,-0.120791), (52270,-0.305139), (52271,-0.277674), (52272,-0.489429), (52273,-0.544643), (52274,-0.298871), (52275,-0.043343), (52276,-0.212363), (52277,-0.234133), (52278,-0.275421), (52279,-0.111858), (52280,-0.412329), (52281,-0.489847), (52282,-0.205984), (52283,0.040257), (52284,-0.110184), (52285,-0.196988), (52286,-0.357642), (52287,-0.355730), (52288,-0.507562), (52289,-0.553953), (52290,-0.330015), (52291,-0.012703), (52292,-0.169650), (52293,-0.233230), (52294,-0.295876), (52295,-0.163903), (52296,-0.395627), (52297,-0.450384), (52298,-0.157230), (52299,0.098762), (52300,-0.051210), (52301,-0.090175), (52302,-0.300997), (52303,-0.330200), (52304,-0.453704), (52305,-0.512637), (52306,-0.255249), (52307,0.016071), (52308,-0.106963), (52309,-0.184938), (52310,-0.241085), (52311,-0.088211), (52312,-0.431417), (52313,-0.493137), (52314,-0.239932), (52315,0.010956), (52316,-0.120907), (52317,-0.165438), (52318,-0.333531), (52319,-0.333010), (52320,-0.488561), (52321,-0.548884), (52322,-0.318440), (52323,-0.025286), (52324,-0.178514), (52325,-0.225838), (52326,-0.312642), (52327,-0.163481), (52328,-0.515047), (52329,-0.181943), (52330,-0.330061), (52331,-0.047126), (52332,-0.220328), (52333,-0.295986), (52334,-0.436672), (52335,-0.417103), (52336,-0.535027), (52337,-0.231660), (52338,-0.373736), (52339,-0.127963), (52340,-0.283977), (52341,-0.264408), (52342,-0.447830), (52343,-0.247573), (52344,-0.439354), (52345,-0.501074), (52346,-0.261801), (52347,0.018811), (52348,-0.146959), (52349,-0.191496), (52350,-0.366552), (52351,-0.408297), (52352,-0.713414), (52353,-0.757019), (52354,-0.544690), (52355,-0.267328), (52356,-0.472114), (52357,-0.472056), (52358,-0.560720), (52359,-0.428747), (52360,-0.860669), (52361,-0.495055), (52362,-0.649209), (52363,-0.382072), (52364,-0.511142), (52365,-0.588191), (52366,-0.693109), (52367,-0.744147), (52368,-0.863004), (52369,-0.558234), (52370,-0.691024), (52371,-0.426673), (52372,-0.571535), (52373,-0.576124), (52374,-0.677793), (52375,-0.564862), (52376,-0.652599), (52377,-0.680411), (52378,-0.445785), (52379,-0.155880), (52380,-0.325827), (52381,-0.404271), (52382,-0.581650), (52383,-0.574629), (52384,-0.744112), (52385,-0.803509), (52386,-0.577711), (52387,-0.297099), (52388,-0.433602), (52389,-0.464201), (52390,-0.529177), (52391,-0.394418), (52392,-0.718113), (52393,-0.472334), (52394,-0.570754), (52395,-0.673813), (52396,-0.402030), (52397,-0.586372), (52398,-0.670859), (52399,-0.795283), (52400,-0.783616), (52401,-0.522515), (52402,-0.544748), (52403,-0.702159), (52404,-0.441985), (52405,-0.501381), (52406,-0.568210), (52407,-0.689391), (52408,-0.645670), (52409,-0.702744), (52410,-0.506670), (52411,-0.222808), (52412,-0.374640), (52413,-0.372728), (52414,-0.579838), (52415,-0.569560), (52416,-0.752976), (52417,-0.806806), (52418,-0.602830), (52419,-0.306426), (52420,-0.471732), (52421,-0.518123), (52422,-0.567301), (52423,-0.407464), (52424,-0.640578), (52425,-0.429646), (52426,-0.441197), (52427,-0.625545), (52428,-0.361658), (52429,-0.544146), (52430,-0.581251), (52431,-0.747015), (52432,-0.746030), (52433,-0.492362), (52434,-0.548972), (52435,-0.758404), (52436,-0.446672), (52437,-0.530689), (52438,-0.586366), (52439,-0.705687), (52440,-0.648961), (52441,-0.687926), (52442,-0.422172), (52443,-0.175010), (52444,-0.335200), (52445,-0.380201), (52446,-0.560367), (52447,-0.554736), (52448,-0.734438), (52449,-0.715802), (52450,-0.496967), (52451,-0.184308), (52452,-0.378875), (52453,-0.472178), (52454,-0.545050), (52455,-0.400999), (52456,-0.429275), (52457,-0.574606), (52458,-0.239186), (52459,-0.386371), (52460,-0.116441), (52461,-0.289644), (52462,-0.383417), (52463,-0.505054), (52464,-0.503606), (52465,-0.621994), (52466,-0.237338), (52467,-0.431905), (52468,-0.160579), (52469,-0.306374), (52470,-0.231533), (52471,-0.417277), (52472,-0.473424), (52473,-0.579270), (52474,-0.320492), (52475,-0.052422), (52476,-0.183815), (52477,-0.259010), (52478,-0.397373), (52479,-0.419143), (52480,-0.685243), (52481,-0.705623), (52482,-0.444059), (52483,-0.139759), (52484,-0.301346), (52485,-0.396973), (52486,-0.459156), (52487,-0.307678), (52488,-0.487380), (52489,-0.629456), (52490,-0.221112), (52491,-0.389662), (52492,-0.101153), (52493,-0.292934), (52494,-0.366733), (52495,-0.526460), (52496,-0.538017), (52497,-0.689385), (52498,-0.348392), (52499,-0.497437), (52500,-0.171772), (52501,-0.360296), (52502,-0.322155), (52503,-0.469340), (52504,-0.549175), (52505,-0.615077), (52506,-0.359086), (52507,-0.083583), (52508,-0.205690), (52509,-0.243722), (52510,-0.453612), (52511,-0.452627), (52512,-0.618860), (52513,-0.688946), (52514,-0.445490), (52515,-0.127258), (52516,-0.327861), (52517,-0.388654), (52518,-0.418320), (52519,-0.264056), (52520,-0.483701), (52521,-0.512910), (52522,-0.292679), (52523,-0.041334), (52524,-0.209891), (52525,-0.229338), (52526,-0.383029), (52527,-0.392263), (52528,-0.527376), (52529,-0.620679), (52530,-0.366548), (52531,-0.066424), (52532,-0.200610), (52533,-0.266512), (52534,-0.342164), (52535,-0.181857), (52536,-0.516705), (52537,-0.623477), (52538,-0.372132), (52539,-0.088270), (52540,-0.222913), (52541,-0.274883), (52542,-0.506608), (52543,-0.499580), (52544,-0.652808), (52545,-0.688053), (52546,-0.450177), (52547,-0.167705), (52548,-0.306067), (52549,-0.366397), (52550,-0.389564), (52551,-0.239939), (52552,-0.489785), (52553,-0.524560), (52554,-0.313158), (52555,-0.028369), (52556,-0.156976), (52557,-0.209410), (52558,-0.383069), (52559,-0.405309), (52560,-0.569683), (52561,-0.635122), (52562,-0.367052), (52563,-0.128712), (52564,-0.276824), (52565,-0.323685), (52566,-0.394227), (52567,-0.243213), (52568,-0.503734), (52569,-0.566387), (52570,-0.310859), (52571,-0.010735), (52572,-0.175115), (52573,-0.269815), (52574,-0.454626), (52575,-0.445276), (52576,-0.590144), (52577,-0.623067), (52578,-0.404695), (52579,-0.145454), (52580,-0.287993), (52581,-0.355292), (52582,-0.401683), (52583,-0.252985), (52584,-0.617094), (52585,-0.268204), (52586,-0.436754), (52587,-0.166361), (52588,-0.332131), (52589,-0.440300), (52590,-0.591204), (52591,-0.591616), (52592,-0.744837), (52593,-0.399661), (52594,-0.511549), (52595,-0.257881), (52596,-0.386024), (52597,-0.392003), (52598,-0.508074), (52599,-0.354730), (52600,-0.556730), (52601,-0.619382), (52602,-0.340160), (52603,-0.065127), (52604,-0.231354), (52605,-0.318158), (52606,-0.499720), (52607,-0.432775), (52608,-0.801529), (52609,-0.881364), (52610,-0.627696), (52611,-0.341974), (52612,-0.509597), (52613,-0.546702), (52614,-0.613531), (52615,-0.461120), (52616,-0.610629), (52617,-0.647734), (52618,-0.417753), (52619,-0.126459), (52620,-0.287119), (52621,-0.350229), (52622,-0.539687), (52623,-0.521050), (52624,-0.696106), (52625,-0.778270), (52626,-0.484652), (52627,-0.223545), (52628,-0.399071), (52629,-0.430597), (52630,-0.470025), (52631,-0.364063), (52632,-0.682649), (52633,-0.708139), (52634,-0.478622), (52635,-0.214271), (52636,-0.383284), (52637,-0.391592), (52638,-0.575940), (52639,-0.531293), (52640,-0.693806), (52641,-0.745770), (52642,-0.517650), (52643,-0.237964), (52644,-0.417203), (52645,-0.436656), (52646,-0.521137), (52647,-0.353398), (52648,-0.462500), (52649,-0.620367), (52650,-0.276587), (52651,-0.396835), (52652,-0.114363), (52653,-0.268987), (52654,-0.364613), (52655,-0.525274), (52656,-0.549837), (52657,-0.676584), (52658,-0.354169), (52659,-0.535730), (52660,-0.278806), (52661,-0.414382), (52662,-0.386453), (52663,-0.522493), (52664,-0.744467), (52665,-0.797364), (52666,-0.557165), (52667,-0.239853), (52668,-0.422811), (52669,-0.447374), (52670,-0.612674), (52671,-0.608440), (52672,-0.769094), (52673,-0.826637), (52674,-0.606406), (52675,-0.315111), (52676,-0.469272), (52677,-0.523559), (52678,-0.597357), (52679,-0.435191), (52680,-0.446279), (52681,-0.597183), (52682,-0.234825), (52683,-0.411277), (52684,-0.157603), (52685,-0.348920), (52686,-0.414823), (52687,-0.559685), (52688,-0.541975), (52689,-0.679874), (52690,-0.353746), (52691,-0.493962), (52692,-0.230538), (52693,-0.413959), (52694,-0.369312), (52695,-0.504418), (52696,-0.706882), (52697,-0.766285), (52698,-0.498215), (52699,-0.208310), (52700,-0.329484), (52701,-0.369376), (52702,-0.581595), (52703,-0.552739), (52704,-0.689242), (52705,-0.782552), (52706,-0.532597), (52707,-0.249198), (52708,-0.437259), (52709,-0.498052), (52710,-0.560235), (52711,-0.394819), (52712,-0.457935), (52713,-0.645996), (52714,-0.283638), (52715,-0.439182), (52716,-0.147424), (52717,-0.283001), (52718,-0.336361), (52719,-0.499808), (52720,-0.505786), (52721,-0.627430), (52722,-0.283180), (52723,-0.507008), (52724,-0.212927), (52725,-0.369405), (52726,-0.380962), (52727,-0.560201), (52728,-0.393388), (52729,-0.471833), (52730,-0.588367), (52731,0.094501), (52732,-0.040611), (52733,-0.119519), (52734,-0.277393), (52735,-0.307992), (52736,-0.335342), (52737,-0.359898), (52738,-0.514522), (52739,0.133969), (52740,-0.021112), (52741,-0.089801), (52742,-0.229096), (52743,-0.034413), (52744,-0.225730), (52745,-0.370592), (52746,-0.415130), (52747,-0.189789), (52748,0.088500), (52749,-0.030821), (52750,-0.101833), (52751,-0.301040), (52752,-0.288910), (52753,-0.451893), (52754,-0.498284), (52755,-0.252506), (52756,0.005809), (52757,-0.157175), (52758,-0.172445), (52759,-0.279687), (52760,-0.367418), (52761,-0.423565), (52762,-0.614419), (52763,0.080522), (52764,-0.082918), (52765,-0.152540), (52766,-0.315054), (52767,-0.309886), (52768,-0.478906), (52769,-0.555028), (52770,-0.679921), (52771,0.016416), (52772,-0.108014), (52773,-0.194818), (52774,-0.330858), (52775,-0.117133), (52776,-0.581572), (52777,-0.590806), (52778,-0.329236), (52779,-0.024472), (52780,-0.216716), (52781,-0.260784), (52782,-0.485545), (52783,-0.450654), (52784,-0.601552), (52785,-0.658168), (52786,-0.386842), (52787,-0.131314), (52788,-0.255281), (52789,-0.327683), (52790,-0.376397), (52791,-0.215627), (52792,-0.347020), (52793,-0.419892), (52794,-0.574047), (52795,0.099529), (52796,-0.065777), (52797,-0.116814), (52798,-0.285371), (52799,-0.328512), (52800,-0.475234), (52801,-0.523948), (52802,-0.683675), (52803,-0.011032), (52804,-0.145682), (52805,-0.202292), (52806,-0.328575), (52807,-0.110204), (52808,-0.342398), (52809,-0.406441), (52810,-0.546200), (52811,0.149211), (52812,0.038713), (52813,-0.034152), (52814,-0.197599), (52815,-0.218906), (52816,-0.403718), (52817,-0.442682), (52818,-0.593587), (52819,0.050728), (52820,-0.119224), (52821,-0.135422), (52822,-0.299332), (52823,-0.072138), (52824,-0.351244), (52825,-0.372551), (52826,-0.528565), (52827,0.125500), (52828,-0.022155), (52829,-0.073192), (52830,-0.257077), (52831,-0.250977), (52832,-0.414887), (52833,-0.497045), (52834,-0.615439), (52835,0.069283), (52836,-0.071866), (52837,-0.127549), (52838,-0.245474), (52839,-0.013634), (52840,-0.426044), (52841,-0.450144), (52842,-0.225737), (52843,0.046980), (52844,-0.066298), (52845,-0.111763), (52846,-0.271027), (52847,-0.297449), (52848,-0.440458), (52849,-0.489172), (52850,-0.263368), (52851,0.021884), (52852,-0.138307), (52853,-0.193527), (52854,-0.280794), (52855,-0.139529), (52856,-0.520826), (52857,-0.597874), (52858,-0.377643), (52859,-0.044082), (52860,-0.199633), (52861,-0.254383), (52862,-0.423403), (52863,-0.427065), (52864,-0.623485), (52865,-0.690321), (52866,-0.477059), (52867,-0.133742), (52868,-0.326450), (52869,-0.344044), (52870,-0.423415), (52871,-0.315593), (52872,-0.589590), (52873,-0.323843), (52874,-0.390672), (52875,-0.599635), (52876,-0.271647), (52877,-0.447173), (52878,-0.509356), (52879,-0.682088), (52880,-0.699682), (52881,-0.389346), (52882,-0.480796), (52883,-0.609866), (52884,-0.364094), (52885,-0.393766), (52886,-0.420646), (52887,-0.591988), (52888,-0.379660), (52889,-0.566794), (52890,-0.264348), (52891,-0.425008), (52892,-0.119781), (52893,-0.272539), (52894,-0.333795), (52895,-0.479127), (52896,-0.532488), (52897,-0.647162), (52898,-0.316851), (52899,-0.473792), (52900,-0.206648), (52901,-0.327359), (52902,-0.329161), (52903,-0.480992), (52904,-0.610069), (52905,-0.393557), (52906,-0.442272), (52907,-0.598286), (52908,-0.284693), (52909,-0.448603), (52910,-0.529834), (52911,-0.670520), (52912,-0.619830), (52913,-0.415397), (52914,-0.417662), (52915,-0.606657), (52916,-0.327441), (52917,-0.394733), (52918,-0.451344), (52919,-0.587846), (52920,-0.485604), (52921,-0.625826), (52922,-0.262065), (52923,-0.427372), (52924,-0.130041), (52925,-0.334358), (52926,-0.416985), (52927,-0.584608), (52928,-0.524169), (52929,-0.657422), (52930,-0.343366), (52931,-0.510989), (52932,-0.234097), (52933,-0.341802), (52934,-0.350567), (52935,-0.495435), (52936,-0.542759), (52937,-0.361545), (52938,-0.374498), (52939,-0.514714), (52940,-0.205305), (52941,-0.386866), (52942,-0.456482), (52943,-0.570693), (52944,-0.590610), (52945,-0.325790), (52946,-0.371717), (52947,-0.524945), (52948,-0.249906), (52949,-0.340893), (52950,-0.393789), (52951,-0.528896), (52952,-0.392283), (52953,-0.544115), (52954,-0.199865), (52955,-0.337764), (52956,-0.081310), (52957,-0.240110), (52958,-0.319481), (52959,-0.479209), (52960,-0.468932), (52961,-0.579423), (52962,-0.241216), (52963,-0.438570), (52964,-0.163531), (52965,-0.335800), (52966,-0.254923), (52967,-0.385389), (52968,-0.275251), (52969,-0.415930), (52970,-0.075864), (52971,-0.256499), (52972,0.031546), (52973,-0.125864), (52974,-0.199656), (52975,-0.375182), (52976,-0.347253), (52977,-0.478183), (52978,-0.164597), (52979,-0.318752), (52980,-0.036743), (52981,-0.203909), (52982,-0.171798), (52983,-0.369621), (52984,-0.327290), (52985,-0.508389), (52986,-0.184114), (52987,-0.331769), (52988,-0.042797), (52989,-0.193696), (52990,-0.261921), (52991,-0.433264), (52992,-0.412768), (52993,-0.612908), (52994,-0.254726), (52995,-0.405631), (52996,-0.161248), (52997,-0.340487), (52998,-0.274938), (52999,-0.415161), (53000,-0.419749), (53001,-0.553465), (53002,-0.193887), (53003,-0.347115), (53004,-0.074398), (53005,-0.251314), (53006,-0.312107), (53007,-0.474627), (53008,-0.447162), (53009,-0.607822), (53010,-0.281224), (53011,-0.410294), (53012,-0.147333), (53013,-0.302421), (53014,-0.263810), (53015,-0.380808), (53016,-0.510811), (53017,-0.565098), (53018,-0.309106), (53019,-0.021061), (53020,-0.179862), (53021,-0.206742), (53022,-0.369725), (53023,-0.358521), (53024,-0.568417), (53025,-0.632460), (53026,-0.356957), (53027,-0.069376), (53028,-0.244901), (53029,-0.290366), (53030,-0.382279), (53031,-0.253093), (53032,-0.404924), (53033,-0.448992), (53034,-0.238523), (53035,0.026297), (53036,-0.209610), (53037,-0.201192), (53038,-0.384144), (53039,-0.312553), (53040,-0.489938), (53041,-0.555841), (53042,-0.276618), (53043,-0.010408), (53044,-0.158063), (53045,-0.205381), (53046,-0.294044), (53047,-0.114690), (53048,-0.505742), (53049,-0.516366), (53050,-0.295672), (53051,-0.003914), (53052,-0.159928), (53053,-0.219788), (53054,-0.408319), (53055,-0.380860), (53056,-0.558702), (53057,-0.587442), (53058,-0.350492), (53059,-0.063380), (53060,-0.210102), (53061,-0.280651), (53062,-0.376277), (53063,-0.221080), (53064,-0.433762), (53065,-0.479690), (53066,-0.247387), (53067,0.011391), (53068,-0.155306), (53069,-0.182185), (53070,-0.373503), (53071,-0.370658), (53072,-0.484869), (53073,-0.538693), (53074,-0.290598), (53075,-0.033210), (53076,-0.163677), (53077,-0.217964), (53078,-0.314060), (53079,-0.156540), (53080,-0.446322), (53081,-0.507578), (53082,-0.241368), (53083,0.007191), (53084,-0.146500), (53085,-0.195678), (53086,-0.423225), (53087,-0.404589), (53088,-0.556883), (53089,-0.603744), (53090,-0.374227), (53091,-0.084786), (53092,-0.253342), (53093,-0.287191), (53094,-0.367495), (53095,-0.204402), (53096,-0.464460), (53097,-0.218688), (53098,-0.248354), (53099,-0.432702), (53100,-0.134445), (53101,-0.301141), (53102,-0.335454), (53103,-0.500760), (53104,-0.498842), (53105,-0.249814), (53106,-0.292492), (53107,-0.468481), (53108,-0.166040), (53109,-0.250052), (53110,-0.292266), (53111,-0.432488), (53112,-0.406883), (53113,-0.461170), (53114,-0.214001), (53115,0.080080), (53116,-0.082903), (53117,-0.132544), (53118,-0.306673), (53119,-0.296866), (53120,-0.175112), (53121,0.063697), (53122,0.036348), (53123,-0.147068), (53124,0.087559), (53125,0.031412), (53126,-0.008943), (53127,-0.159384), (53128,-0.134248), (53129,0.121286), (53130,0.081858), (53131,-0.090411), (53132,0.148861), (53133,-0.046169), (53134,-0.061909), (53135,-0.208631), (53136,-0.202074), (53137,0.018157), (53138,-0.024984), (53139,-0.162883), (53140,0.142813), (53141,0.088057), (53142,0.059781), (53143,-0.145006), (53144,-0.108254), (53145,0.130555), (53146,0.093450), (53147,-0.064887), (53148,0.231517), (53149,0.051815), (53150,-0.030343), (53151,-0.171028), (53152,-0.162148), (53153,0.094777), (53154,0.046526), (53155,-0.114598), (53156,0.178557), (53157,0.095466), (53158,0.037002), (53159,-0.116225), (53160,0.216872), (53161,0.101734), (53162,-0.021300), (53163,-0.055618), (53164,-0.253436), (53165,-0.003017), (53166,-0.133947), (53167,-0.182198), (53168,0.072867), (53169,0.057133), (53170,-0.084943), (53171,-0.141096), (53172,-0.187487), (53173,0.054109), (53174,-0.104692), (53175,-0.187313), (53176,-0.153348), (53177,0.103107), (53178,0.026985), (53179,-0.106268), (53180,0.182704), (53181,-0.002571), (53182,-0.011805), (53183,-0.191507), (53184,-0.229539), (53185,0.053396), (53186,-0.007397), (53187,-0.163411), (53188,0.121848), (53189,0.074524), (53190,-0.006701), (53191,-0.166435), (53192,-0.023773), (53193,0.305141), (53194,0.126366), (53195,0.038635), (53196,-0.100654), (53197,0.168343), (53198,-0.006250), (53199,-0.037775), (53200,-0.186827), (53201,0.206659), (53202,0.100350), (53203,0.056275), (53204,-0.091373), (53205,0.236615), (53206,0.070382), (53207,-0.011776), (53208,-0.117622), (53209,0.148125), (53210,0.068754), (53211,-0.090980), (53212,0.198462), (53213,0.036874), (53214,-0.000694), (53215,-0.160428), (53216,-0.158510), (53217,0.116060), (53218,0.077101), (53219,-0.091455), (53220,0.174762), (53221,0.093994), (53222,0.026232), (53223,-0.133032), (53224,0.043073), (53225,0.345977), (53226,0.237808), (53227,0.137066), (53228,0.010782), (53229,0.242622), (53230,0.094040), (53231,0.015132), (53232,-0.129266), (53233,0.295803), (53234,0.137002), (53235,0.081782), (53236,-0.064476), (53237,0.291382), (53238,0.178104), (53239,0.101519), (53240,-0.021978), (53241,0.262347), (53242,0.199231), (53243,0.045077), (53244,0.300605), (53245,0.129269), (53246,0.090767), (53247,-0.106587), (53248,-0.085157), (53249,0.147609), (53250,0.130479), (53251,-0.022749), (53252,0.264833), (53253,0.172456), (53254,0.068000), (53255,-0.051784), (53256,-0.061945), (53257,0.276262), (53258,0.112816), (53259,0.071534), (53260,-0.084017), (53261,0.191949), (53262,0.018290), (53263,0.001160), (53264,-0.164610), (53265,0.261855), (53266,0.114200), (53267,0.091034), (53268,-0.067304), (53269,0.325718), (53270,0.131151), (53271,0.044347), (53272,0.103396), (53273,-0.028930), (53274,0.283266), (53275,0.144904), (53276,0.438985), (53277,0.262532), (53278,0.230543), (53279,0.091248), (53280,0.025352), (53281,-0.118120), (53282,0.227983), (53283,0.076151), (53284,0.355367), (53285,0.217931), (53286,0.231928), (53287,0.051756), (53288,0.010475), (53289,0.272972), (53290,0.210319), (53291,0.100754), (53292,0.353965), (53293,0.196091), (53294,0.106964), (53295,-0.077384), (53296,-0.057351), (53297,0.199104), (53298,0.148999), (53299,-0.057647), (53300,0.237367), (53301,0.171928), (53302,0.141793), (53303,-0.086682), (53304,-0.090806), (53305,0.131278), (53306,0.098819), (53307,-0.064621), (53308,0.233173), (53309,0.077628), (53310,-0.035656), (53311,-0.166123), (53312,-0.177674), (53313,0.054630), (53314,0.038889), (53315,-0.099473), (53316,0.154665), (53317,0.058569), (53318,0.038188), (53319,-0.148013), (53320,-0.107549), (53321,0.146126), (53322,0.118313), (53323,-0.043280), (53324,0.231296), (53325,0.072495), (53326,0.033074), (53327,-0.156854), (53328,-0.155400), (53329,0.096879), (53330,0.015184), (53331,-0.101350), (53332,0.218742), (53333,0.084099), (53334,0.051640), (53335,-0.074180), (53336,0.056866), (53337,-0.117727), (53338,0.267856), (53339,0.114628), (53340,0.404533), (53341,0.260134), (53342,0.182616), (53343,0.040541), (53344,0.056854), (53345,-0.079186), (53346,0.272490), (53347,0.110903), (53348,0.378973), (53349,0.170937), (53350,0.238346), (53351,0.097660), (53352,0.310922), (53353,0.131220), (53354,0.055098), (53355,-0.072582), (53356,0.201994), (53357,0.047370), (53358,-0.022709), (53359,-0.150389), (53360,0.263071), (53361,0.116806), (53362,0.033259), (53363,-0.142730), (53364,0.230780), (53365,0.102173), (53366,0.053922), (53367,-0.098842), (53368,0.048929), (53369,0.270080), (53370,0.239481), (53371,0.049560), (53372,0.329709), (53373,0.149544), (53374,0.118475), (53375,-0.077946), (53376,-0.161500), (53377,0.133508), (53378,0.000724), (53379,0.179610), (53380,0.047747), (53381,0.047805), (53382,-0.112386), (53383,0.137106), (53384,-0.079759), (53385,0.253338), (53386,0.075496), (53387,0.096919), (53388,-0.069315), (53389,-0.156119), (53390,-0.316309), (53391,-0.025015), (53392,-0.150835), (53393,0.208737), (53394,0.065728), (53395,0.182842), (53396,-0.008475), (53397,0.060330), (53398,-0.107763), (53399,0.152411), (53400,-0.122049), (53401,0.134412), (53402,0.100557), (53403,-0.095401), (53404,-0.028925), (53405,-0.206304), (53406,-0.273133), (53407,-0.429148), (53408,-0.161078), (53409,0.075409), (53410,0.020652), (53411,-0.113991), (53412,-0.022895), (53413,-0.111558), (53414,-0.118933), (53415,-0.242430), (53416,-0.024992), (53417,0.246798), (53418,0.215266), (53419,0.054612), (53420,0.030512), (53421,-0.164982), (53422,-0.174216), (53423,-0.324188), (53424,-0.054728), (53425,0.239817), (53426,0.131648), (53427,-0.014147), (53428,0.100174), (53429,0.033345), (53430,-0.049740), (53431,-0.202504), (53432,-0.063562), (53433,0.165491), (53434,0.114454), (53435,-0.071754), (53436,-0.054044), (53437,-0.223527), (53438,-0.267138), (53439,-0.438474), (53440,-0.125815), (53441,0.101379), (53442,0.039196), (53443,-0.106136), (53444,0.042562), (53445,-0.017304), (53446,-0.043721), (53447,-0.191376), (53448,0.035355), (53449,0.272768), (53450,0.239382), (53451,0.087551), (53452,0.106187), (53453,-0.099532), (53454,-0.153356), (53455,-0.301004), (53456,-0.089602), (53457,0.204479), (53458,0.152509), (53459,0.007183), (53460,0.162844), (53461,0.066748), (53462,0.043118), (53463,-0.101751), (53464,-0.067786), (53465,0.143153), (53466,0.069818), (53467,-0.096409), (53468,-0.087992), (53469,-0.227751), (53470,-0.285757), (53471,-0.448734), (53472,-0.143971), (53473,0.078577), (53474,0.047515), (53475,-0.127541), (53476,0.008608), (53477,-0.042893), (53478,-0.090211), (53479,-0.268523), (53480,0.019986), (53481,0.270404), (53482,0.217044), (53483,0.082864), (53484,0.085239), (53485,-0.091677), (53486,-0.132495), (53487,-0.323806), (53488,-0.041804), (53489,0.193756), (53490,0.152931), (53491,0.008069), (53492,0.135396), (53493,0.061597), (53494,0.016603), (53495,-0.115260), (53496,0.242922), (53497,0.093877), (53498,0.413505), (53499,0.297904), (53500,0.292853), (53501,0.187470), (53502,0.083478), (53503,-0.061390), (53504,0.190888), (53505,0.046489), (53506,0.370764), (53507,0.165978), (53508,0.346722), (53509,0.161911), (53510,0.207955), (53511,0.109072), (53512,0.190876), (53513,0.052513), (53514,0.383758), (53515,0.208702), (53516,0.212473), (53517,0.085720), (53518,-0.004798), (53519,-0.185426), (53520,0.129556), (53521,-0.033891), (53522,0.337760), (53523,0.158058), (53524,0.287714), (53525,0.140522), (53526,0.194926), (53527,0.042161), (53528,0.097961), (53529,0.016730), (53530,0.220236), (53531,0.204502), (53532,0.049414), (53533,0.032284), (53534,-0.117688), (53535,0.182893), (53536,0.002264), (53537,-0.071071), (53538,0.182604), (53539,0.340124), (53540,0.218017), (53541,0.144682), (53542,0.041623), (53543,0.348709), (53544,-0.066494), (53545,0.255457), (53546,0.112918), (53547,0.127835), (53548,-0.032819), (53549,-0.096398), (53550,-0.232438), (53551,0.042596), (53552,-0.103663), (53553,0.215502), (53554,0.092932), (53555,0.198894), (53556,0.069360), (53557,0.135372), (53558,-0.038757), (53559,0.194943), (53560,0.063550), (53561,0.047346), (53562,0.323775), (53563,0.332193), (53564,0.163173), (53565,0.068943), (53566,-0.061993), (53567,0.236734), (53568,0.032881), (53569,0.000885), (53570,0.198355), (53571,0.322432), (53572,0.188246), (53573,0.146037), (53574,0.068519), (53575,0.361211), (53576,0.123914), (53577,0.100741), (53578,0.339087), (53579,0.333102), (53580,0.206355), (53581,0.120478), (53582,-0.078736), (53583,0.231144), (53584,0.038900), (53585,-0.007498), (53586,0.220166), (53587,0.373040), (53588,0.199374), (53589,0.152056), (53590,0.103806), (53591,0.382558), (53592,0.116921), (53593,0.031050), (53594,0.240592), (53595,0.284776), (53596,0.136658), (53597,0.094913), (53598,-0.114983), (53599,0.214865), (53600,0.080679), (53601,0.042184), (53602,0.288889), (53603,0.381382), (53604,0.246269), (53605,0.216134), (53606,0.123757), (53607,0.393217), (53608,0.063022), (53609,0.383114), (53610,0.231746), (53611,0.259675), (53612,0.107374), (53613,0.008497), (53614,-0.148913), (53615,0.135418), (53616,0.013311), (53617,0.345482), (53618,0.204333), (53619,0.315404), (53620,0.193760), (53621,0.218903), (53622,0.070321), (53623,0.321666), (53624,-0.002029), (53625,0.292052), (53626,0.153226), (53627,0.146315), (53628,0.070193), (53629,-0.010568), (53630,-0.174941), (53631,0.075477), (53632,-0.202233), (53633,0.070014), (53634,0.015263), (53635,-0.149110), (53636,0.001904), (53637,-0.028231), (53638,-0.102493), (53639,-0.262221), (53640,0.020709), (53641,0.280883), (53642,0.221023), (53643,0.013913), (53644,0.006075), (53645,-0.150865), (53646,-0.198190), (53647,-0.381605), (53648,-0.060123), (53649,0.178687), (53650,0.127186), (53651,-0.065521), (53652,0.110114), (53653,0.023310), (53654,-0.038879), (53655,-0.182815), (53656,-0.406179), (53657,0.259501), (53658,0.128571), (53659,0.087746), (53660,-0.103102), (53661,-0.098397), (53662,-0.266027), (53663,-0.339356), (53664,-0.497230), (53665,0.168444), (53666,0.030082), (53667,-0.029778), (53668,-0.210407), (53669,0.048371), (53670,-0.091852), (53671,-0.085757), (53672,-0.318408), (53673,0.355631), (53674,0.175923), (53675,0.121636), (53676,-0.012080), (53677,-0.093775), (53678,-0.222382), (53679,-0.266919), (53680,-0.387630), (53681,0.292446), (53682,0.140151), (53683,0.066816), (53684,-0.103594), (53685,0.083187), (53686,-0.035201), (53687,-0.062550), (53688,-0.439200), (53689,0.255277), (53690,0.077435), (53691,0.018502), (53692,-0.142159), (53693,-0.105871), (53694,-0.264208), (53695,-0.361231), (53696,-0.513062), (53697,0.160507), (53698,0.008213), (53699,-0.041898), (53700,-0.229496), (53701,0.032538), (53702,-0.124403), (53703,-0.187519), (53704,-0.291511), (53705,0.370919), (53706,0.260421), (53707,0.154575), (53708,-0.003298), (53709,0.006515), (53710,-0.189442), (53711,-0.235370), (53712,-0.380238), (53713,0.323062), (53714,0.170304), (53715,0.108578), (53716,-0.051149), (53717,0.209951), (53718,0.010744), (53719,-0.047262), (53720,-0.437845), (53721,0.230622), (53722,0.082503), (53723,0.049581), (53724,-0.089714), (53725,-0.131923), (53726,-0.317204), (53727,-0.367308), (53728,-0.491738), (53729,0.147931), (53730,-0.028985), (53731,-0.068876), (53732,-0.182624), (53733,0.057112), (53734,-0.111438), (53735,-0.140184), (53736,-0.336605), (53737,0.354153), (53738,0.213005), (53739,0.172650), (53740,-0.007516), (53741,-0.027896), (53742,-0.200635), (53743,-0.252136), (53744,-0.401644), (53745,0.240342), (53746,0.109876), (53747,0.039327), (53748,-0.098566), (53749,0.131414), (53750,-0.009271), (53751,-0.076564), (53752,-0.101590), (53753,0.188308), (53754,0.395997), (53755,0.328698), (53756,0.155966), (53757,0.221051), (53758,0.062250), (53759,-0.012938), (53760,-0.168489), (53761,0.114910), (53762,0.344890), (53763,0.321724), (53764,0.174069), (53765,0.322766), (53766,0.236426), (53767,0.229515), (53768,-0.142953), (53769,0.152524), (53770,0.385755), (53771,0.364911), (53772,0.211220), (53773,0.241466), (53774,0.050618), (53775,0.014446), (53776,-0.132746), (53777,0.125569), (53778,0.378780), (53779,0.304981), (53780,0.166156), (53781,0.325066), (53782,0.243372), (53783,0.195584), (53784,0.249060), (53785,0.111625), (53786,0.456338), (53787,0.264557), (53788,0.293882), (53789,0.115570), (53790,0.036662), (53791,-0.122602), (53792,0.164510), (53793,-0.025411), (53794,0.339277), (53795,0.208347), (53796,0.354715), (53797,0.210779), (53798,0.222916), (53799,0.073402), (53800,0.042339), (53801,0.319238), (53802,0.258909), (53803,0.107077), (53804,0.165194), (53805,-0.030764), (53806,-0.074375), (53807,-0.237352), (53808,0.037218), (53809,0.277424), (53810,0.237995), (53811,0.066189), (53812,0.226496), (53813,0.125297), (53814,0.085405), (53815,-0.095693), (53816,0.236014), (53817,0.055385), (53818,0.408921), (53819,0.239901), (53820,0.255751), (53821,0.102524), (53822,0.019433), (53823,-0.150050), (53824,0.113844), (53825,-0.009190), (53826,0.321584), (53827,0.192044), (53828,0.306835), (53829,0.174509), (53830,0.210797), (53831,0.086836), (53832,0.308457), (53833,0.182167), (53834,0.493436), (53835,0.309552), (53836,0.315182), (53837,0.151272), (53838,0.051463), (53839,-0.071571), (53840,0.182567), (53841,0.046064), (53842,0.399600), (53843,0.261237), (53844,0.351407), (53845,0.229300), (53846,0.244686), (53847,0.077990), (53848,0.273130), (53849,0.119439), (53850,0.485987), (53851,0.336942), (53852,0.323988), (53853,0.200027), (53854,0.096968), (53855,-0.060443), (53856,0.230389), (53857,0.084130), (53858,0.433490), (53859,0.266793), (53860,0.407588), (53861,0.259007), (53862,0.257668), (53863,0.173657), (53864,0.181605), (53865,0.399049), (53866,0.328037), (53867,0.178059), (53868,0.254297), (53869,0.069949), (53870,0.054215), (53871,-0.136639), (53872,0.176490), (53873,0.394391), (53874,0.348927), (53875,0.173408), (53876,0.317923), (53877,0.224149), (53878,0.160570), (53879,0.031500), (53880,0.043630), (53881,0.295445), (53882,0.238372), (53883,0.104186), (53884,0.108890), (53885,-0.030869), (53886,-0.114886), (53887,-0.253712), (53888,-0.137531), (53889,0.103131), (53890,0.049771), (53891,-0.120639), (53892,0.017840), (53893,-0.031807), (53894,-0.082381), (53895,-0.235609), (53896,-0.077156), (53897,0.150965), (53898,0.105037), (53899,-0.071415), (53900,-0.038377), (53901,-0.199964), (53902,-0.261220), (53903,-0.441386), (53904,-0.179821), (53905,0.094291), (53906,0.083661), (53907,-0.106724), (53908,0.050797), (53909,-0.036934), (53910,-0.080545), (53911,-0.242595), (53912,-0.247184), (53913,0.036215), (53914,0.267592), (53915,0.186824), (53916,0.051718), (53917,0.075927), (53918,-0.111671), (53919,-0.137167), (53920,-0.297821), (53921,-0.020928), (53922,0.232746), (53923,0.180776), (53924,0.052169), (53925,0.203190), (53926,0.108954), (53927,0.048161), (53928,-0.274608), (53929,0.417083), (53930,0.233661), (53931,0.130139), (53932,-0.034235), (53933,-0.027677), (53934,-0.181832), (53935,-0.185030), (53936,-0.313173), (53937,0.331606), (53938,0.170482), (53939,0.113872), (53940,-0.063507), (53941,0.212922), (53942,0.069450), (53943,-0.002489), (53944,-0.422802), (53945,0.223367), (53946,0.078035), (53947,0.036290), (53948,-0.143875), (53949,-0.187486), (53950,-0.323525), (53951,-0.365270), (53952,-0.518498), (53953,0.149969), (53954,-0.003259), (53955,-0.047797), (53956,-0.209384), (53957,0.015957), (53958,-0.147954), (53959,-0.171590), (53960,-0.350359), (53961,0.323681), (53962,0.167666), (53963,0.065534), (53964,-0.038458), (53965,-0.076490), (53966,-0.274770), (53967,-0.309089), (53968,-0.431190), (53969,0.228911), (53970,0.022265), (53971,0.006531), (53972,-0.168062), (53973,0.091186), (53974,-0.030458), (53975,-0.101470), (53976,-0.254698), (53977,0.042639), (53978,0.223848), (53979,0.190462), (53980,0.066965), (53981,0.101856), (53982,-0.086205), (53983,-0.141425), (53984,-0.270032), (53985,-0.011254), (53986,0.203867), (53987,0.176048), (53988,0.021431), (53989,0.170592), (53990,0.081001), (53991,0.080126), (53992,-0.138129), (53993,0.118795), (53994,0.366427), (53995,0.274051), (53996,0.144511), (53997,0.120418), (53998,-0.060217), (53999,-0.070379), (54000,-0.224533), (54001,0.066762), (54002,0.293956), (54003,0.261960), (54004,0.098050), (54005,0.244425), (54006,0.144615), (54007,0.140027), (54008,-0.064296), (54009,0.221895), (54010,0.459308), (54011,0.412448), (54012,0.221137), (54013,0.244882), (54014,0.083759), (54015,0.035045), (54016,-0.154413), (54017,0.101115), (54018,0.341314), (54019,0.296313), (54020,0.137513), (54021,0.282491), (54022,0.219381), (54023,0.175776), (54024,-0.153498), (54025,0.120614), (54026,0.376606), (54027,0.313953), (54028,0.175127), (54029,0.197946), (54030,0.002916), (54031,-0.042085), (54032,-0.207385), (54033,0.064398), (54034,0.273477), (54035,0.241488), (54036,0.105912), (54037,0.269005), (54038,0.181737), (54039,0.118621), (54040,0.086626), (54041,-0.040585), (54042,0.281361), (54043,0.123957), (54044,0.154209), (54045,0.009340), (54046,-0.074214), (54047,-0.207930), (54048,-0.009534), (54049,-0.152079), (54050,0.181488), (54051,0.039406), (54052,0.227584), (54053,0.115702), (54054,0.112040), (54055,-0.032822), (54056,0.222706), (54057,0.059259), (54058,0.360310), (54059,0.208472), (54060,0.186239), (54061,0.052986), (54062,-0.046361), (54063,-0.132238), (54064,0.095420), (54065,-0.034577), (54066,0.304556), (54067,0.156438), (54068,0.302349), (54069,0.152841), (54070,0.192842), (54071,0.026609), (54072,0.207354), (54073,0.037408), (54074,0.326379), (54075,0.188480), (54076,0.242883), (54077,0.074796), (54078,-0.023623), (54079,-0.179637), (54080,0.075428), (54081,-0.088946), (54082,0.304076), (54083,0.191261), (54084,0.333453), (54085,0.147245), (54086,0.151016), (54087,0.041921), (54088,0.233348), (54089,0.096375), (54090,0.391389), (54091,0.267422), (54092,0.236823), (54093,0.084529), (54094,-0.014354), (54095,-0.153643), (54096,0.136255), (54097,-0.003498), (54098,0.308235), (54099,0.175446), (54100,0.325070), (54101,0.162086), (54102,0.184906), (54103,0.048866), (54104,0.136250), (54105,0.013216), (54106,0.338417), (54107,0.141527), (54108,0.175028), (54109,0.046885), (54110,-0.012981), (54111,-0.173172), (54112,0.091648), (54113,-0.068085), (54114,0.255726), (54115,0.096926), (54116,0.243764), (54117,0.101682), (54118,0.099880), (54119,-0.025477), (54120,0.112075), (54121,0.382468), (54122,0.320742), (54123,0.148936), (54124,0.197303), (54125,-0.011660), (54126,-0.036223), (54127,-0.234040), (54128,0.025201), (54129,0.319752), (54130,0.284507), (54131,0.115487), (54132,0.231668), (54133,0.169015), (54134,0.121691), (54135,-0.028281), (54136,0.002434), (54137,0.239847), (54138,0.169299), (54139,0.059734), (54140,0.075120), (54141,-0.136635), (54142,-0.179777), (54143,-0.368765), (54144,-0.031484), (54145,-0.171707), (54146,0.177183), (54147,0.002127), (54148,0.153611), (54149,0.002706), (54150,0.053860), (54151,-0.106801), (54152,-0.235877), (54153,0.060997), (54154,0.266356), (54155,0.186985), (54156,0.022611), (54157,0.049144), (54158,-0.140314), (54159,-0.197851), (54160,-0.327854), (54161,-0.037023), (54162,0.224542), (54163,0.186046), (54164,0.027709), (54165,0.172694), (54166,0.060342), (54167,0.054358), (54168,-0.306031), (54169,-0.045394), (54170,0.166008), (54171,0.118221), (54172,0.005406), (54173,0.037511), (54174,-0.167739), (54175,-0.226208), (54176,-0.414270), (54177,-0.137840), (54178,0.133016), (54179,0.102417), (54180,-0.104692), (54181,0.036109), (54182,-0.028397), (54183,-0.033918), (54184,-0.346461), (54185,0.303884), (54186,0.157625), (54187,0.110771), (54188,-0.076364), (54189,-0.108359), (54190,-0.254154), (54191,-0.294973), (54192,-0.487680), (54193,0.216083), (54194,0.095836), (54195,0.012288), (54196,-0.158128), (54197,0.092754), (54198,-0.058144), (54199,-0.099896), (54200,-0.281458), (54201,0.018666), (54202,0.217989), (54203,0.153947), (54204,-0.035974), (54205,-0.012692), (54206,-0.187284), (54207,-0.262016), (54208,-0.411061), (54209,-0.109084), (54210,0.102788), (54211,0.065220), (54212,-0.077789), (54213,0.089950), (54214,0.020335), (54215,-0.021880), (54216,-0.200655), (54217,0.047446), (54218,0.294145), (54219,0.242181), (54220,0.097776), (54221,0.110840), (54222,-0.065612), (54223,-0.090632), (54224,-0.261048), (54225,-0.072408), (54226,0.182657), (54227,0.164600), (54228,-0.008133), (54229,0.122444), (54230,0.075589), (54231,0.038484), (54232,-0.357671), (54233,-0.059408), (54234,0.159890), (54235,0.094451), (54236,-0.103829), (54237,-0.061505), (54238,-0.262108), (54239,-0.304786), (54240,-0.427357), (54241,-0.228497), (54242,0.023318), (54243,-0.046304), (54244,-0.187916), (54245,-0.050834), (54246,-0.119523), (54247,-0.173347), (54248,-0.362341), (54249,-0.034347), (54250,0.211425), (54251,0.142737), (54252,-0.044398), (54253,-0.013683), (54254,-0.200354), (54255,-0.232813), (54256,-0.420875), (54257,-0.130976), (54258,0.154746), (54259,0.083270), (54260,-0.049983), (54261,0.103824), (54262,0.032349), (54263,-0.012652), (54264,-0.219292), (54265,0.087332), (54266,0.314989), (54267,0.255123), (54268,0.087036), (54269,0.115891), (54270,-0.084712), (54271,-0.167803), (54272,-0.258320), (54273,0.018573), (54274,0.290826), (54275,0.217491), (54276,0.060087), (54277,0.198095), (54278,0.138236), (54279,0.083015), (54280,-0.241613), (54281,0.065943), (54282,0.308466), (54283,0.258355), (54284,0.098165), (54285,0.075925), (54286,-0.078230), (54287,-0.111152), (54288,-0.261130), (54289,0.011586), (54290,0.253182), (54291,0.179847), (54292,0.035448), (54293,0.185999), (54294,0.124280), (54295,0.089498), (54296,0.330161), (54297,0.137916), (54298,0.046003), (54299,0.264374), (54300,0.267682), (54301,0.112601), (54302,0.060631), (54303,-0.107926), (54304,0.192661), (54305,0.026891), (54306,-0.005561), (54307,0.245321), (54308,0.378690), (54309,0.215243), (54310,0.155840), (54311,0.092267), (54312,0.074667), (54313,-0.041861), (54314,0.287060), (54315,0.105962), (54316,0.094868), (54317,-0.049068), (54318,-0.105215), (54319,-0.273771), (54320,0.043071), (54321,-0.136631), (54322,0.219698), (54323,0.050215), (54324,0.210985), (54325,0.048465), (54326,0.075930), (54327,-0.068005), (54328,0.073253), (54329,-0.046994), (54330,0.295866), (54331,0.168649), (54332,0.172420), (54333,-0.007745), (54334,-0.087117), (54335,-0.232912), (54336,0.054200), (54337,-0.042823), (54338,0.254978), (54339,0.123584), (54340,0.260203), (54341,0.083751), (54342,0.114929), (54343,-0.035512), (54344,0.116899), (54345,-0.075809), (54346,0.327896), (54347,0.196496), (54348,0.155214), (54349,0.014529), (54350,-0.086207), (54351,-0.238972), (54352,0.056969), (54353,-0.086040), (54354,0.282361), (54355,0.118451), (54356,0.294087), (54357,0.115311), (54358,0.163215), (54359,0.020669), (54360,0.346341), (54361,0.197289), (54362,0.161117), (54363,0.372519), (54364,0.380937), (54365,0.223533), (54366,0.185037), (54367,-0.013713), (54368,0.291984), (54369,0.108099), (54370,0.051489), (54371,0.279146), (54372,0.454318), (54373,0.307133), (54374,0.266315), (54375,0.201802), (54376,0.133577), (54377,0.412799), (54378,0.344573), (54379,0.154189), (54380,0.149137), (54381,-0.019882), (54382,-0.060700), (54383,-0.222757), (54384,0.074117), (54385,0.289232), (54386,0.229835), (54387,0.063139), (54388,0.277327), (54389,0.155683), (54390,0.107896), (54391,-0.099671), (54392,0.165143), (54393,0.017025), (54394,0.388682), (54395,0.221053), (54396,0.196959), (54397,0.079035), (54398,-0.028207), (54399,-0.171216), (54400,-0.353704), (54401,-0.068916), (54402,0.157352), (54403,0.109101), (54404,-0.047377), (54405,0.071591), (54406,0.027523), (54407,-0.029557), (54408,-0.278006), (54409,0.015148), (54410,0.254884), (54411,0.211743), (54412,0.014389), (54413,0.046964), (54414,-0.122989), (54415,-0.173093), (54416,-0.359764), (54417,-0.049891), (54418,0.187985), (54419,0.124412), (54420,0.008341), (54421,0.189086), (54422,0.080454), (54423,0.000619), (54424,-0.310540), (54425,-0.061975), (54426,0.173578), (54427,0.152271), (54428,-0.013035), (54429,-0.015300), (54430,-0.191753), (54431,-0.215383), (54432,-0.426205), (54433,-0.132587), (54434,0.135946), (54435,0.077476), (54436,-0.074825), (54437,0.085488), (54438,-0.036619), (54439,-0.089053), (54440,-0.231128), (54441,0.034156), (54442,0.274355), (54443,0.200093), (54444,0.044079), (54445,0.056679), (54446,-0.132779), (54447,-0.125758), (54448,-0.354695), (54449,-0.063864), (54450,0.180518), (54451,0.194508), (54452,0.009697), (54453,0.187655), (54454,0.133832), (54455,0.048418), (54456,-0.344025), (54457,-0.026249), (54458,0.229742), (54459,0.203326), (54460,0.055207), (54461,-0.039492), (54462,-0.157886), (54463,-0.237721), (54464,-0.368188), (54465,-0.058308), (54466,0.175385), (54467,0.133177), (54468,-0.051171), (54469,0.104026), (54470,0.029294), (54471,-0.028706), (54472,-0.174037), (54473,0.092173), (54474,0.308684), (54475,0.287378), (54476,0.091414), (54477,0.146280), (54478,-0.077084), (54479,-0.085386), (54480,-0.215389), (54481,0.044785), (54482,0.297990), (54483,0.241380), (54484,0.068647), (54485,0.172749), (54486,0.106847), (54487,0.081357), (54488,-0.355211), (54489,-0.085281), (54490,0.126584), (54491,0.121996), (54492,-0.041914), (54493,-0.036283), (54494,-0.193224), (54495,-0.256804), (54496,-0.401209), (54497,-0.172618), (54498,0.094988), (54499,0.023050), (54500,-0.146903), (54501,0.009691), (54502,-0.076650), (54503,-0.144406), (54504,-0.206595), (54505,-0.338915), (54506,0.365775), (54507,0.218590), (54508,0.174985), (54509,0.006429), (54510,0.021352), (54511,-0.156496), (54512,-0.214966), (54513,-0.384913), (54514,0.290054), (54515,0.134039), (54516,0.076503), (54517,-0.075329), (54518,0.156511), (54519,-0.021801), (54520,-0.216368), (54521,0.043343), (54522,0.271463), (54523,0.233432), (54524,0.076954), (54525,0.100700), (54526,-0.079465), (54527,-0.155124), (54528,-0.295339), (54529,-0.017520), (54530,0.249160), (54531,0.224597), (54532,0.047682), (54533,0.184300), (54534,0.173213), (54535,0.125889), (54536,-0.102122), (54537,-0.296226), (54538,0.383856), (54539,0.256639), (54540,0.234399), (54541,0.069099), (54542,0.065438), (54543,-0.082217), (54544,-0.188990), (54545,-0.306451), (54546,0.334608), (54547,0.157693), (54548,0.137313), (54549,0.022175), (54550,0.231254), (54551,0.071057), (54552,0.252265), (54553,0.120408), (54554,0.055902), (54555,0.331868), (54556,0.382552), (54557,0.202850), (54558,0.129051), (54559,-0.033462), (54560,0.256436), (54561,0.059545), (54562,0.045208), (54563,0.248244), (54564,0.377900), (54565,0.218630), (54566,0.194073), (54567,0.117489), (54568,-0.214103), (54569,0.098557), (54570,0.349438), (54571,0.277036), (54572,0.077359), (54573,0.068125), (54574,-0.117150), (54575,-0.116165), (54576,-0.288898), (54577,-0.046375), (54578,0.190574), (54579,0.114453), (54580,-0.007655), (54581,0.167517), (54582,0.088146), (54583,0.074266), (54584,0.146784), (54585,-0.001328), (54586,0.344775), (54587,0.245429), (54588,0.264065), (54589,0.095509), (54590,-0.027525), (54591,-0.155205), (54592,0.111012), (54593,-0.068227), (54594,0.248152), (54595,0.120935), (54596,0.212965), (54597,0.107113), (54598,0.130859), (54599,-0.005181), (54600,-0.145866), (54601,0.087833), (54602,0.367976), (54603,0.315085), (54604,0.140956), (54605,0.118253), (54606,-0.027542), (54607,-0.037703), (54608,-0.207186), (54609,0.048805), (54610,0.304796), (54611,0.294172), (54612,0.083349), (54613,0.235297), (54614,0.165675), (54615,0.134149), (54616,0.396177), (54617,0.222981), (54618,0.136177), (54619,0.377772), (54620,0.401982), (54621,0.239931), (54622,0.184248), (54623,0.009186), (54624,0.301413), (54625,0.131467), (54626,0.085533), (54627,0.291825), (54628,0.461425), (54629,0.271040), (54630,0.237654), (54631,0.166179), (54632,-0.083197), (54633,0.172795), (54634,0.398592), (54635,0.390291), (54636,0.239386), (54637,0.253377), (54638,0.021189), (54639,0.016138), (54640,-0.123158), (54641,0.135157), (54642,0.355851), (54643,0.322465), (54644,0.147873), (54645,0.283095), (54646,0.222766), (54647,0.199599), (54648,-0.126883), (54649,0.155589), (54650,0.369314), (54651,0.348465), (54652,0.183164), (54653,0.209233), (54654,0.000728), (54655,-0.060992), (54656,-0.258346), (54657,0.033412), (54658,0.247607), (54659,0.200283), (54660,0.025227), (54661,0.197143), (54662,0.144716), (54663,0.051406), (54664,-0.203080), (54665,0.097971), (54666,0.364645), (54667,0.296889), (54668,0.131119), (54669,0.152078), (54670,0.019752), (54671,-0.086094), (54672,-0.286697), (54673,0.046864), (54674,0.287063), (54675,0.248105), (54676,0.059580), (54677,0.215704), (54678,0.134936), (54679,0.099691), (54680,-0.207280), (54681,0.056608), (54682,0.254078), (54683,0.251349), (54684,0.127382), (54685,0.139049), (54686,-0.056445), (54687,-0.127920), (54688,-0.302049), (54689,0.016189), (54690,0.239201), (54691,0.181200), (54692,-0.005934), (54693,0.130215), (54694,0.070355), (54695,0.038359), (54696,-0.086065), (54697,-0.224897), (54698,0.439857), (54699,0.283842), (54700,0.213294), (54701,0.097693), (54702,0.052692), (54703,-0.083811), (54704,-0.128812), (54705,-0.262065), (54706,0.426839), (54707,0.256423), (54708,0.178912), (54709,0.000600), (54710,0.259847), (54711,0.111266), (54712,-0.110709), (54713,-0.224914), (54714,0.449125), (54715,0.315872), (54716,0.250433), (54717,0.080024), (54718,0.062893), (54719,-0.113096), (54720,-0.176675), (54721,-0.314111), (54722,0.381300), (54723,0.222963), (54724,0.106428), (54725,-0.029611), (54726,0.192010), (54727,0.062007), (54728,-0.051272), (54729,-0.211462), (54730,0.495551), (54731,0.360908), (54732,0.314047), (54733,0.135278), (54734,0.117678), (54735,-0.009532), (54736,-0.083331), (54737,-0.241668), (54738,0.462565), (54739,0.331635), (54740,0.265733), (54741,0.119005), (54742,0.384288), (54743,0.238500), (54744,-0.083342), (54745,-0.277910), (54746,0.372905), (54747,0.241975), (54748,0.155171), (54749,-0.002233), (54750,-0.030515), (54751,-0.147507), (54752,-0.231987), (54753,-0.376856), (54754,0.285105), (54755,0.135596), (54756,0.075267), (54757,-0.103039), (54758,0.109290), (54759,0.007157), (54760,-0.066178), (54761,-0.182242), (54762,0.453244), (54763,0.333460), (54764,0.281496), (54765,0.141274), (54766,0.109741), (54767,-0.049523), (54768,-0.057824), (54769,-0.248678), (54770,0.437440), (54771,0.247982), (54772,0.201128), (54773,0.050223), (54774,0.256979), (54775,0.161353), (54776,0.027630), (54777,-0.108873), (54778,0.573526), (54779,0.420298), (54780,0.346036), (54781,0.219753), (54782,0.229097), (54783,0.052181), (54784,-0.031367), (54785,-0.255201), (54786,0.399333), (54787,0.302310), (54788,0.222006), (54789,0.097582), (54790,0.341495), (54791,0.196632), (54792,-0.057389), (54793,-0.196215), (54794,0.492220), (54795,0.354320), (54796,0.250798), (54797,0.105003), (54798,0.112493), (54799,-0.027265), (54800,-0.085272), (54801,-0.217129), (54802,0.453191), (54803,0.285105), (54804,0.212233), (54805,0.067834), (54806,0.294565), (54807,0.134368), (54808,0.024803), (54809,0.310061), (54810,0.157297), (54811,0.509442), (54812,0.330667), (54813,0.341871), (54814,0.195612), (54815,0.148295), (54816,-0.018865), (54817,0.281252), (54818,0.137317), (54819,0.458805), (54820,0.311150), (54821,0.448232), (54822,0.287109), (54823,0.288563), (54824,-0.141506), (54825,0.147466), (54826,0.423902), (54827,0.379827), (54828,0.169468), (54829,0.178349), (54830,0.005153), (54831,-0.050994), (54832,-0.205149), (54833,0.090792), (54834,0.310090), (54835,0.268802), (54836,0.129050), (54837,0.316764), (54838,0.211375), (54839,0.138973), (54840,-0.117835), (54841,0.155345), (54842,0.390898), (54843,0.336611), (54844,0.188029), (54845,0.182045), (54846,-0.004620), (54847,-0.037542), (54848,-0.182874), (54849,0.136754), (54850,0.359302), (54851,0.315698), (54852,0.131813), (54853,0.235921), (54854,0.200212), (54855,0.112012), (54856,-0.170807), (54857,0.142785), (54858,0.354651), (54859,0.353312), (54860,0.197761), (54861,0.208502), (54862,0.044592), (54863,-0.027810), (54864,-0.195434), (54865,0.093068), (54866,0.349066), (54867,0.312888), (54868,0.180568), (54869,0.320900), (54870,0.222023), (54871,0.201174), (54872,0.102761), (54873,0.335527), (54874,0.212030), (54875,0.559060), (54876,0.416521), (54877,0.432371), (54878,0.273570), (54879,0.195589), (54880,0.042831), (54881,0.288140), (54882,0.126553), (54883,0.491704), (54884,0.343122), (54885,0.482528), (54886,0.331623), (54887,0.381380), (54888,0.013089), (54889,0.274196), (54890,0.538546), (54891,0.462895), (54892,0.316166), (54893,0.335736), (54894,0.122590), (54895,0.073406), (54896,-0.095144), (54897,0.217516), (54898,0.454002), (54899,0.441518), (54900,0.246487), (54901,0.416543), (54902,0.323240), (54903,0.248045), (54904,-0.045457), (54905,0.203109), (54906,0.484648), (54907,0.403417), (54908,0.285492), (54909,0.293909), (54910,0.120244), (54911,0.059451), (54912,-0.247057), (54913,0.021014), (54914,0.225446), (54915,0.168836), (54916,-0.002507), (54917,0.173592), (54918,0.076106), (54919,0.030178), (54920,-0.243812), (54921,0.030758), (54922,0.280249), (54923,0.264046), (54924,0.109891), (54925,0.128991), (54926,-0.007975), (54927,-0.063195), (54928,-0.233605), (54929,0.027959), (54930,0.272342), (54931,0.212945), (54932,0.057394), (54933,0.187507), (54934,0.103026), (54935,0.095652), (54936,-0.160693), (54937,-0.265612), (54938,0.411677), (54939,0.281217), (54940,0.123806), (54941,0.012851), (54942,0.027768), (54943,-0.129636), (54944,-0.216904), (54945,-0.358986), (54946,0.310408), (54947,0.134425), (54948,0.108936), (54949,-0.055444), (54950,0.188011), (54951,0.005523), (54952,-0.074318), (54953,-0.229863), (54954,0.440921), (54955,0.302558), (54956,0.191603), (54957,0.056490), (54958,0.041220), (54959,-0.118508), (54960,-0.213671), (54961,-0.305121), (54962,0.397716), (54963,0.208258), (54964,0.173939), (54965,0.024431), (54966,0.257668), (54967,0.142060), (54968,-0.098956), (54969,-0.281445), (54970,0.415819), (54971,0.229148), (54972,0.203658), (54973,0.063906), (54974,0.012868), (54975,-0.133390), (54976,-0.176068), (54977,-0.364599), (54978,0.347993), (54979,0.176187), (54980,0.094956), (54981,-0.046656), (54982,0.187507), (54983,0.039852), (54984,-0.028837), (54985,-0.232690), (54986,0.472007), (54987,0.339680), (54988,0.270528), (54989,0.098722), (54990,0.133614), (54991,-0.000566), (54992,-0.117564), (54993,-0.268932), (54994,0.442264), (54995,0.269068), (54996,0.223141), (54997,0.012781), (54998,0.249725), (54999,0.129014), (55000,-0.151482), (55001,-0.329325), (55002,0.361897), (55003,0.192414), (55004,0.153918), (55005,-0.011851), (55006,-0.043841), (55007,-0.179417), (55008,-0.231850), (55009,-0.384615), (55010,0.296394), (55011,0.132947), (55012,0.104671), (55013,-0.049947), (55014,0.168888), (55015,-0.001991), (55016,-0.066497), (55017,-0.207646), (55018,0.463600), (55019,0.321061), (55020,0.262591), (55021,0.097748), (55022,0.087587), (55023,-0.061921), (55024,-0.128750), (55025,-0.255967), (55026,0.386952), (55027,0.237907), (55028,0.177114), (55029,0.053610), (55030,0.238075), (55031,0.067665), (55032,0.160152), (55033,0.012033), (55034,0.297292), (55035,0.576977), (55036,0.526867), (55037,0.349024), (55038,0.352796), (55039,0.149406), (55040,0.053773), (55041,-0.075297), (55042,0.239222), (55043,0.468275), (55044,0.415842), (55045,0.273766), (55046,0.444292), (55047,0.344013), (55048,0.138300), (55049,-0.027000), (55050,0.244783), (55051,0.465477), (55052,0.392142), (55053,0.235665), (55054,0.292854), (55055,0.075062), (55056,0.031921), (55057,-0.119447), (55058,0.156982), (55059,0.347020), (55060,0.351254), (55061,0.192923), (55062,0.344871), (55063,0.254811), (55064,-0.007571), (55065,0.257250), (55066,0.086834), (55067,0.421328), (55068,0.246735), (55069,0.287206), (55070,0.169282), (55071,0.094087), (55072,-0.044276), (55073,0.215898), (55074,0.061281), (55075,0.399951), (55076,0.242084), (55077,0.395884), (55078,0.236157), (55079,0.256183), (55080,-0.179452), (55081,0.125775), (55082,0.359938), (55083,0.292182), (55084,0.119443), (55085,0.143652), (55086,-0.005856), (55087,-0.066185), (55088,-0.227309), (55089,0.069565), (55090,0.252633), (55091,0.250831), (55092,0.083201), (55093,0.222607), (55094,0.149741), (55095,0.094058), (55096,-0.009934), (55097,0.254423), (55098,0.103518), (55099,0.487247), (55100,0.320551), (55101,0.330358), (55102,0.173881), (55103,0.103338), (55104,-0.036884), (55105,0.209358), (55106,0.044515), (55107,0.388301), (55108,0.267590), (55109,0.374015), (55110,0.211959), (55111,0.253826), (55112,-0.002989), (55113,0.244650), (55114,0.097458), (55115,0.489547), (55116,0.312168), (55117,0.300147), (55118,0.127878), (55119,0.100992), (55120,-0.046193), (55121,0.240455), (55122,0.139719), (55123,0.438446), (55124,0.280572), (55125,0.457604), (55126,0.289511), (55127,0.285386), (55128,0.034620), (55129,0.299904), (55130,0.161542), (55131,0.485347), (55132,0.331192), (55133,0.319635), (55134,0.173840), (55135,0.100511), (55136,-0.095453), (55137,0.238578), (55138,0.109508), (55139,0.418448), (55140,0.274976), (55141,0.395339), (55142,0.240722), (55143,0.284436), (55144,-0.016962), (55145,0.213482), (55146,0.465760), (55147,0.424942), (55148,0.270324), (55149,0.286174), (55150,0.093467), (55151,0.028028), (55152,-0.153071), (55153,0.140083), (55154,0.400258), (55155,0.333428), (55156,0.183451), (55157,0.317746), (55158,0.275075), (55159,0.228677), (55160,-0.086189), (55161,0.212538), (55162,0.444378), (55163,0.389622), (55164,0.214566), (55165,0.235988), (55166,0.039098), (55167,0.001066), (55168,-0.366292), (55169,-0.079643), (55170,0.164276), (55171,0.103019), (55172,-0.007473), (55173,0.148188), (55174,0.064171), (55175,0.035431), (55176,-0.245071), (55177,0.005353), (55178,0.229291), (55179,0.222386), (55180,0.068226), (55181,0.076180), (55182,-0.108632), (55183,-0.161992), (55184,-0.349590), (55185,-0.033675), (55186,0.192123), (55187,0.107642), (55188,0.028734), (55189,0.184401), (55190,0.076226), (55191,0.013579), (55192,0.028496), (55193,-0.125658), (55194,0.126620), (55195,0.370069), (55196,0.346903), (55197,0.199718), (55198,0.211385), (55199,0.016817), (55200,-0.065340), (55201,-0.196270), (55202,0.097348), (55203,0.377027), (55204,0.258176), (55205,0.106344), (55206,0.262005), (55207,0.135258), (55208,-0.072315), (55209,-0.183276), (55210,0.485653), (55211,0.333359), (55212,0.301827), (55213,0.137916), (55214,0.096172), (55215,-0.024076), (55216,-0.087655), (55217,-0.240420), (55218,0.402036), (55219,0.245095), (55220,0.226105), (55221,0.081706), (55222,0.294035), (55223,0.106437), (55224,-0.202863), (55225,-0.355621), (55226,0.300767), (55227,0.211640), (55228,0.129482), (55229,-0.018173), (55230,-0.053882), (55231,-0.204323), (55232,-0.245605), (55233,-0.419734), (55234,0.271957), (55235,0.123839), (55236,0.081161), (55237,-0.100864), (55238,0.161170), (55239,-0.069164), (55240,-0.123914), (55241,-0.279465), (55242,0.403397), (55243,0.235774), (55244,0.176377), (55245,0.064489), (55246,0.069656), (55247,-0.114228), (55248,-0.214501), (55249,-0.331499), (55250,0.364369), (55251,0.173984), (55252,0.136879), (55253,0.017565), (55254,0.203419), (55255,0.051588), (55256,-0.048691), (55257,-0.172652), (55258,0.104241), (55259,0.356519), (55260,0.304555), (55261,0.126713), (55262,0.160208), (55263,-0.008812), (55264,-0.093293), (55265,-0.262312), (55266,0.018300), (55267,0.270578), (55268,0.199566), (55269,0.060277), (55270,0.254954), (55271,0.149108), (55272,0.069274), (55273,-0.065376), (55274,0.224992), (55275,0.470301), (55276,0.402076), (55277,0.260464), (55278,0.287923), (55279,0.091965), (55280,0.041391), (55281,-0.139237), (55282,0.128833), (55283,0.401079), (55284,0.338433), (55285,0.187992), (55286,0.306495), (55287,0.237807), (55288,0.166331), (55289,-0.000365), (55290,0.251913), (55291,0.497222), (55292,0.464300), (55293,0.289244), (55294,0.316703), (55295,0.125392), (55296,-0.249869), (55297,0.041895), (55298,-0.094144), (55299,0.233844), (55300,0.057855), (55301,0.204230), (55302,0.041246), (55303,0.086363), (55304,-0.172305), (55305,-0.299521), (55306,-0.009154), (55307,0.257520), (55308,0.240860), (55309,0.069980), (55310,0.099762), (55311,-0.092012), (55312,-0.166274), (55313,-0.283735), (55314,-0.047255), (55315,0.216175), (55316,0.149809), (55317,-0.011314), (55318,0.144810), (55319,0.070548), (55320,-0.259654), (55321,0.000990), (55322,-0.139232), (55323,0.168781), (55324,0.017413), (55325,-0.003430), (55326,-0.128324), (55327,-0.195616), (55328,-0.367422), (55329,-0.077054), (55330,-0.227959), (55331,0.123717), (55332,-0.055522), (55333,0.099675), (55334,-0.034041), (55335,0.015716), (55336,-0.202076), (55337,0.072963), (55338,-0.096983), (55339,0.224506), (55340,0.075454), (55341,0.128004), (55342,-0.015938), (55343,-0.134789), (55344,-0.280121), (55345,0.008388), (55346,-0.132298), (55347,0.227280), (55348,0.062907), (55349,0.172118), (55350,0.023073), (55351,0.079799), (55352,-0.200233), (55353,0.061331), (55354,-0.077495), (55355,0.249566), (55356,0.112594), (55357,0.129840), (55358,-0.037320), (55359,-0.111582), (55360,-0.272705), (55361,-0.000922), (55362,-0.142998), (55363,0.234689), (55364,0.051737), (55365,0.202752), (55366,0.072755), (55367,0.094178), (55368,-0.117578), (55369,0.162571), (55370,-0.016204), (55371,0.293675), (55372,0.154843), (55373,0.163260), (55374,0.016538), (55375,-0.054937), (55376,-0.206768), (55377,0.043650), (55378,-0.071951), (55379,0.277871), (55380,0.108852), (55381,0.274268), (55382,0.130333), (55383,0.154078), (55384,-0.230468), (55385,0.080338), (55386,-0.113766), (55387,0.231410), (55388,0.043349), (55389,0.075918), (55390,-0.068018), (55391,-0.161791), (55392,-0.278319), (55393,-0.006072), (55394,-0.178342), (55395,0.155689), (55396,-0.014264), (55397,0.123288), (55398,0.002571), (55399,0.012848), (55400,-0.237454), (55401,0.071022), (55402,0.264779), (55403,0.171006), (55404,0.008022), (55405,0.050816), (55406,-0.180914), (55407,-0.210117), (55408,-0.332688), (55409,-0.034887), (55410,0.174192), (55411,0.100394), (55412,-0.058407), (55413,0.076815), (55414,0.005340), (55415,-0.049410), (55416,-0.474370), (55417,-0.139412), (55418,0.106360), (55419,0.067402), (55420,-0.108587), (55421,-0.084841), (55422,-0.283585), (55423,-0.297466), (55424,-0.510611), (55425,-0.201665), (55426,0.002304), (55427,-0.097968), (55428,-0.221929), (55429,-0.092743), (55430,-0.170261), (55431,-0.270070), (55432,-0.647647), (55433,0.058909), (55434,-0.117080), (55435,-0.149076), (55436,-0.314839), (55437,-0.293880), (55438,-0.463832), (55439,-0.502791), (55440,-0.647189), (55441,0.001302), (55442,-0.191405), (55443,-0.235480), (55444,-0.417041), (55445,-0.157794), (55446,-0.295230), (55447,-0.343944), (55448,-0.296973), (55449,-0.463207), (55450,0.174603), (55451,0.048319), (55452,0.001458), (55453,-0.157806), (55454,-0.168430), (55455,-0.304006), (55456,-0.365726), (55457,-0.527313), (55458,0.117460), (55459,-0.082681), (55460,-0.107244), (55461,-0.247459), (55462,0.007135), (55463,-0.177213), (55464,-0.516700), (55465,-0.242124), (55466,0.023623), (55467,-0.199742), (55468,-0.242883), (55469,-0.415153), (55470,-0.380261), (55471,-0.539062), (55472,-0.530644), (55473,-0.282079), (55474,-0.050245), (55475,-0.186285), (55476,-0.259614), (55477,-0.294395), (55478,-0.190294), (55479,-0.333302), (55480,-0.433112), (55481,-0.586339), (55482,0.114181), (55483,-0.014432), (55484,-0.091944), (55485,-0.281865), (55486,-0.256259), (55487,-0.420170), (55488,-0.476780), (55489,-0.591454), (55490,0.041246), (55491,-0.066466), (55492,-0.159306), (55493,-0.289309), (55494,-0.081157), (55495,-0.205118), (55496,-0.415014), (55497,-0.179461), (55498,0.119267), (55499,-0.054399), (55500,-0.118905), (55501,-0.337160), (55502,-0.298549), (55503,-0.460600), (55504,-0.486559), (55505,-0.306277), (55506,-0.007550), (55507,-0.145913), (55508,-0.209492), (55509,-0.257280), (55510,-0.091394), (55511,-0.245085), (55512,-0.295195), (55513,-0.436807), (55514,0.251627), (55515,0.084931), (55516,-0.001410), (55517,-0.159277), (55518,-0.170371), (55519,-0.349147), (55520,-0.454992), (55521,-0.565947), (55522,0.115518), (55523,-0.019125), (55524,-0.088740), (55525,-0.269839), (55526,-0.050078), (55527,-0.132235), (55528,-0.221362), (55529,-0.357402), (55530,0.355191), (55531,0.170379), (55532,0.136061), (55533,-0.040855), (55534,-0.036614), (55535,-0.210280), (55536,-0.275719), (55537,-0.397357), (55538,0.277146), (55539,0.086762), (55540,0.027359), (55541,-0.099852), (55542,0.092039), (55543,-0.044464), (55544,-0.249714), (55545,-0.394119), (55546,0.315224), (55547,0.178252), (55548,0.084021), (55549,-0.065957), (55550,-0.090519), (55551,-0.241887), (55552,-0.340764), (55553,-0.528832), (55554,0.163786), (55555,-0.019166), (55556,-0.036759), (55557,-0.150507), (55558,0.035347), (55559,-0.137849), (55560,-0.334276), (55561,-0.499113), (55562,0.207437), (55563,0.027272), (55564,-0.052563), (55565,-0.183493), (55566,-0.189941), (55567,-0.288823), (55568,-0.374694), (55569,-0.528849), (55570,0.117320), (55571,-0.016396), (55572,-0.065580), (55573,-0.221594), (55574,0.008856), (55575,-0.146695), (55576,-0.451349), (55577,-0.155408), (55578,0.097797), (55579,0.063021), (55580,-0.088347), (55581,-0.024194), (55582,-0.230371), (55583,-0.297663), (55584,-0.462043), (55585,-0.164706), (55586,0.073170), (55587,-0.004804), (55588,-0.156179), (55589,-0.024200), (55590,-0.109614), (55591,-0.137426), (55592,-0.351968), (55593,-0.055095), (55594,0.182782), (55595,0.108983), (55596,-0.025666), (55597,0.020378), (55598,-0.165824), (55599,-0.207575), (55600,-0.358016), (55601,-0.070898), (55602,0.191129), (55603,0.139629), (55604,-0.088382), (55605,0.082144), (55606,0.010668), (55607,-0.025040), (55608,-0.379856), (55609,-0.144297), (55610,0.095903), (55611,0.056938), (55612,-0.105576), (55613,-0.090653), (55614,-0.290799), (55615,-0.329294), (55616,-0.530824), (55617,-0.213055), (55618,0.001596), (55619,-0.009028), (55620,-0.158536), (55621,-0.018204), (55622,-0.056236), (55623,-0.120279), (55624,-0.407744), (55625,-0.096012), (55626,0.129323), (55627,0.093151), (55628,-0.078655), (55629,-0.074884), (55630,-0.269915), (55631,-0.321415), (55632,-0.472784), (55633,-0.166624), (55634,0.077289), (55635,0.034611), (55636,-0.129762), (55637,0.031014), (55638,-0.012127), (55639,-0.079426), (55640,-0.332052), (55641,-0.065378), (55642,0.191546), (55643,0.146545), (55644,-0.023864), (55645,-0.016843), (55646,-0.236958), (55647,-0.287995), (55648,-0.415206), (55649,-0.142026), (55650,0.096777), (55651,0.016015), (55652,-0.125134), (55653,0.025418), (55654,-0.021437), (55655,-0.065048), (55656,-0.489074), (55657,0.240243), (55658,0.092589), (55659,0.010431), (55660,-0.121432), (55661,-0.124161), (55662,-0.275992), (55663,-0.352113), (55664,-0.496982), (55665,0.164515), (55666,0.007575), (55667,-0.069937), (55668,-0.220842), (55669,0.055588), (55670,-0.128291), (55671,-0.166792), (55672,-0.338135), (55673,-0.060309), (55674,0.186860), (55675,0.146505), (55676,-0.043880), (55677,-0.067046), (55678,-0.249535), (55679,-0.254593), (55680,-0.532766), (55681,-0.239148), (55682,0.016843), (55683,-0.058808), (55684,-0.216682), (55685,-0.074491), (55686,-0.170117), (55687,-0.245775), (55688,-0.482146), (55689,-0.150901), (55690,0.073969), (55691,0.017359), (55692,-0.126113), (55693,-0.115372), (55694,-0.312263), (55695,-0.354477), (55696,-0.508168), (55697,-0.208045), (55698,0.020539), (55699,-0.045363), (55700,-0.188835), (55701,-0.046637), (55702,-0.113936), (55703,-0.183088), (55704,-0.428751), (55705,-0.131414), (55706,0.075342), (55707,0.018732), (55708,-0.118240), (55709,-0.122828), (55710,-0.345730), (55711,-0.348458), (55712,-0.502613), (55713,-0.227110), (55714,0.034454), (55715,-0.026802), (55716,-0.185603), (55717,-0.011357), (55718,-0.067504), (55719,-0.133407), (55720,-0.495192), (55721,-0.222476), (55722,0.067423), (55723,-0.059324), (55724,-0.140555), (55725,-0.304002), (55726,-0.319736), (55727,-0.500371), (55728,-0.529111), (55729,-0.298197), (55730,-0.016658), (55731,-0.126223), (55732,-0.186553), (55733,-0.266851), (55734,-0.136275), (55735,-0.277887), (55736,-0.461302), (55737,-0.205774), (55738,0.026529), (55739,-0.068634), (55740,-0.207460), (55741,-0.172105), (55742,-0.342984), (55743,-0.416313), (55744,-0.608094), (55745,-0.301007), (55746,-0.033864), (55747,-0.051927), (55748,-0.207472), (55749,-0.056921), (55750,-0.115854), (55751,-0.191975), (55752,-0.254622), (55753,-0.419465), (55754,0.221594), (55755,0.100884), (55756,-0.002176), (55757,-0.153544), (55758,-0.186002), (55759,-0.301604), (55760,-0.368433), (55761,-0.518411), (55762,0.174207), (55763,-0.022214), (55764,-0.032845), (55765,-0.199541), (55766,0.011398), (55767,-0.110246), (55768,-0.459953), (55769,-0.169122), (55770,0.064115), (55771,-0.025012), (55772,-0.167557), (55773,-0.122910), (55774,-0.305862), (55775,-0.350400), (55776,-0.495725), (55777,-0.243916), (55778,0.019977), (55779,-0.045925), (55780,-0.204263), (55781,-0.078789), (55782,-0.155374), (55783,-0.196662), (55784,-0.199854), (55785,-0.404177), (55786,0.301916), (55787,0.143115), (55788,0.061421), (55789,-0.087630), (55790,-0.078743), (55791,-0.217106), (55792,-0.282545), (55793,-0.425090), (55794,0.213183), (55795,0.065534), (55796,-0.004551), (55797,-0.138268), (55798,0.071738), (55799,-0.091239), (55800,-0.392173), (55801,-0.111561), (55802,0.121206), (55803,0.066449), (55804,-0.056585), (55805,-0.083465), (55806,-0.264100), (55807,-0.349507), (55808,-0.437244), (55809,-0.124578), (55810,0.097969), (55811,0.030207), (55812,-0.103973), (55813,0.028933), (55814,-0.010495), (55815,-0.056886), (55816,-0.244021), (55817,-0.417687), (55818,0.239628), (55819,0.078041), (55820,0.039546), (55821,-0.122505), (55822,-0.128953), (55823,-0.284967), (55824,-0.354582), (55825,-0.506414), (55826,0.160656), (55827,0.038086), (55828,-0.038962), (55829,-0.178252), (55830,0.097715), (55831,-0.037398), (55832,-0.332760), (55833,-0.094420), (55834,0.146713), (55835,0.085456), (55836,-0.079850), (55837,0.005210), (55838,-0.199113), (55839,-0.258510), (55840,-0.408018), (55841,-0.130192), (55842,0.085386), (55843,0.039459), (55844,-0.108660), (55845,0.031679), (55846,-0.059771), (55847,-0.113595), (55848,-0.305376), (55849,-0.074932), (55850,0.231228), (55851,0.181587), (55852,0.020463), (55853,0.013552), (55854,-0.138279), (55855,-0.173988), (55856,-0.350440), (55857,-0.060079), (55858,0.168048), (55859,0.103073), (55860,-0.041790), (55861,0.114804), (55862,0.054011), (55863,0.048953), (55864,-0.348129), (55865,-0.049865), (55866,0.171756), (55867,0.143474), (55868,-0.034832), (55869,-0.026415), (55870,-0.199154), (55871,-0.210705), (55872,-0.412242), (55873,-0.133019), (55874,0.123899), (55875,0.063106), (55876,-0.116596), (55877,0.020956), (55878,-0.042624), (55879,-0.075546), (55880,-0.344896), (55881,-0.056858), (55882,0.186134), (55883,0.105367), (55884,-0.060403), (55885,0.013511), (55886,-0.198708), (55887,-0.285048), (55888,-0.394607), (55889,-0.128397), (55890,0.129918), (55891,0.051010), (55892,-0.115223), (55893,0.051589), (55894,-0.011527), (55895,-0.084856), (55896,-0.344457), (55897,-0.045729), (55898,0.220487), (55899,0.135537), (55900,-0.010258), (55901,0.022317), (55902,-0.156922), (55903,-0.230257), (55904,-0.384412), (55905,-0.120524), (55906,0.111786), (55907,0.044950), (55908,-0.076224), (55909,0.053425), (55910,-0.016654), (55911,-0.066301), (55912,-0.429939), (55913,0.271038), (55914,0.094122), (55915,0.035652), (55916,-0.118966), (55917,-0.137956), (55918,-0.294896), (55919,-0.360799), (55920,-0.486156), (55921,0.196706), (55922,0.082965), (55923,-0.018241), (55924,-0.151494), (55925,0.115186), (55926,-0.043615), (55927,-0.105334), (55928,-0.272501), (55929,-0.006754), (55930,0.245525), (55931,0.202853), (55932,0.056125), (55933,0.046427), (55934,-0.139774), (55935,-0.165264), (55936,-0.583254), (55937,0.076847), (55938,-0.078234), (55939,-0.138564), (55940,-0.295505), (55941,-0.064128), (55942,-0.225252), (55943,-0.256321), (55944,-0.470393), (55945,-0.211146), (55946,0.072717), (55947,-0.098626), (55948,-0.165925), (55949,-0.349340), (55950,-0.310729), (55951,-0.450488), (55952,-0.535896), (55953,-0.331926), (55954,-0.034595), (55955,-0.226840), (55956,-0.267658), (55957,-0.309403), (55958,-0.170461), (55959,-0.323688), (55960,-0.482952), (55961,-0.251582), (55962,0.033677), (55963,-0.114442), (55964,-0.150150), (55965,-0.325670), (55966,-0.338623), (55967,-0.467694), (55968,-0.536382), (55969,-0.311048), (55970,-0.041118), (55971,-0.218034), (55972,-0.223549), (55973,-0.309426), (55974,-0.116602), (55975,-0.299554), (55976,-0.423058), (55977,-0.144299), (55978,0.122838), (55979,-0.029457), (55980,-0.064239), (55981,-0.277848), (55982,-0.239237), (55983,-0.424981), (55984,-0.474159), (55985,-0.211661), (55986,0.060122), (55987,-0.101465), (55988,-0.159008), (55989,-0.228161), (55990,-0.060885), (55991,-0.261488), (55992,-0.570318), (55993,-0.342198), (55994,-0.025819), (55995,-0.195765), (55996,-0.255631), (55997,-0.424651), (55998,-0.390686), (55999,-0.534158), (56000,-0.636291), (56001,-0.393298), (56002,-0.108973), (56003,-0.246872), (56004,-0.283977), (56005,-0.372635), (56006,-0.211401), (56007,-0.327003), (56008,-0.406837), (56009,-0.184289), (56010,0.074488), (56011,-0.080129), (56012,-0.136740), (56013,-0.266743), (56014,-0.282477), (56015,-0.435241), (56016,-0.469090), (56017,-0.240969), (56018,0.032210), (56019,-0.111725), (56020,-0.186450), (56021,-0.271864), (56022,-0.117594), (56023,-0.260602), (56024,-0.465382), (56025,-0.268382), (56026,0.050783), (56027,-0.101981), (56028,-0.174383), (56029,-0.355482), (56030,-0.367502), (56031,-0.489140), (56032,-0.516489), (56033,-0.296728), (56034,-0.049096), (56035,-0.203250), (56036,-0.228740), (56037,-0.299752), (56038,-0.144091), (56039,-0.326117), (56040,-0.386903), (56041,-0.152746), (56042,0.154347), (56043,-0.019319), (56044,-0.098227), (56045,-0.282112), (56046,-0.249537), (56047,-0.419490), (56048,-0.461235), (56049,-0.197811), (56050,0.078619), (56051,-0.052775), (56052,-0.154907), (56053,-0.229169), (56054,-0.085117), (56055,-0.242058), (56056,-0.163041), (56057,-0.271673), (56058,0.357771), (56059,0.226841), (56060,0.117739), (56061,-0.034555), (56062,0.021708), (56063,-0.124088), (56064,-0.220184), (56065,-0.396636), (56066,0.319206), (56067,0.174344), (56068,0.114478), (56069,-0.041530), (56070,0.196810), (56071,0.043582), (56072,-0.146339), (56073,-0.303743), (56074,0.340566), (56075,0.218458), (56076,0.127941), (56077,-0.041078), (56078,-0.060068), (56079,-0.246270), (56080,-0.257828), (56081,-0.418951), (56082,0.274130), (56083,0.132981), (56084,0.048963), (56085,-0.091716), (56086,0.125259), (56087,-0.024256), (56088,-0.299179), (56089,-0.012061), (56090,0.225352), (56091,0.152017), (56092,0.035953), (56093,0.027645), (56094,-0.143698), (56095,-0.237928), (56096,-0.353066), (56097,-0.084532), (56098,0.175172), (56099,0.106489), (56100,-0.035593), (56101,0.097313), (56102,0.067177), (56103,0.011494), (56104,-0.425538), (56105,0.267080), (56106,0.085982), (56107,-0.007792), (56108,-0.115960), (56109,-0.130304), (56110,-0.297464), (56111,-0.368939), (56112,-0.467822), (56113,0.219692), (56114,0.051599), (56115,-0.027772), (56116,-0.183786), (56117,0.024366), (56118,-0.120039), (56119,-0.176649), (56120,-0.265313), (56121,0.012050), (56122,0.270828), (56123,0.245808), (56124,0.083751), (56125,0.061511), (56126,-0.112148), (56127,-0.161796), (56128,-0.357290), (56129,-0.053453), (56130,0.181637), (56131,0.134783), (56132,-0.067681), (56133,0.087517), (56134,0.005359), (56135,-0.056367), (56136,-0.312242), (56137,-0.005619), (56138,0.226221), (56139,0.198408), (56140,0.047040), (56141,0.080072), (56142,-0.121458), (56143,-0.146484), (56144,-0.282993), (56145,-0.036288), (56146,0.156072), (56147,0.133832), (56148,-0.027755), (56149,0.147881), (56150,0.081052), (56151,0.041160), (56152,-0.247702), (56153,0.060781), (56154,0.263361), (56155,0.212787), (56156,0.058632), (56157,0.099097), (56158,-0.069923), (56159,-0.141398), (56160,-0.271865), (56161,0.011071), (56162,0.233155), (56163,0.143101), (56164,-0.012913), (56165,0.158076), (56166,0.056413), (56167,0.046716), (56168,-0.312746), (56169,0.322734), (56170,0.172762), (56171,0.129621), (56172,-0.001773), (56173,-0.041664), (56174,-0.180027), (56175,-0.234783), (56176,-0.382432), (56177,0.260481), (56178,0.147203), (56179,0.079447), (56180,-0.078891), (56181,0.155273), (56182,0.014124), (56183,-0.058748), (56184,-0.482774), (56185,0.233068), (56186,0.072877), (56187,0.000932), (56188,-0.144393), (56189,-0.168029), (56190,-0.324507), (56191,-0.365788), (56192,-0.424722), (56193,-0.589559), (56194,0.071932), (56195,-0.058064), (56196,-0.146728), (56197,-0.315284), (56198,-0.082511), (56199,-0.193473), (56200,-0.349487), (56201,-0.515714), (56202,0.154606), (56203,-0.026492), (56204,-0.068701), (56205,-0.220069), (56206,-0.198646), (56207,-0.409468), (56208,-0.417313), (56209,-0.569607), (56210,0.086317), (56211,-0.032077), (56212,-0.115625), (56213,-0.269316), (56214,-0.025867), (56215,-0.191167), (56216,-0.434506), (56217,-0.511555), (56218,-0.268105), (56219,0.002751), (56220,-0.114247), (56221,-0.164814), (56222,-0.338480), (56223,-0.326349), (56224,-0.502332), (56225,-0.532468), (56226,-0.291805), (56227,-0.027448), (56228,-0.164421), (56229,-0.245652), (56230,-0.344065), (56231,-0.181898), (56232,-0.334199), (56233,-0.384773), (56234,-0.133421), (56235,0.122106), (56236,-0.031585), (56237,-0.050105), (56238,-0.247922), (56239,-0.210707), (56240,-0.388556), (56241,-0.479536), (56242,-0.237941), (56243,0.020374), (56244,-0.138890), (56245,-0.210365), (56246,-0.264189), (56247,-0.114101), (56248,-0.428974), (56249,-0.480475), (56250,-0.217514), (56251,0.032441), (56252,-0.088740), (56253,-0.100754), (56254,-0.273957), (56255,-0.307342), (56256,-0.471252), (56257,-0.488383), (56258,-0.237037), (56259,0.064946), (56260,-0.095714), (56261,-0.138392), (56262,-0.214977), (56263,-0.093224), (56264,-0.296613), (56265,-0.333719), (56266,-0.100482), (56267,0.168978), (56268,0.011111), (56269,-0.057578), (56270,-0.183862), (56271,-0.202389), (56272,-0.348647), (56273,-0.377856), (56274,-0.168771), (56275,0.124377), (56276,-0.060435), (56277,-0.121691), (56278,-0.234506), (56279,-0.058407), (56280,-0.454563), (56281,-0.557158), (56282,-0.296521), (56283,-0.011726), (56284,-0.179355), (56285,-0.226673), (56286,-0.396626), (56287,-0.363588), (56288,-0.508456), (56289,-0.552987), (56290,-0.327190), (56291,-0.030316), (56292,-0.171935), (56293,-0.239227), (56294,-0.285618), (56295,-0.132744), (56296,-0.359828), (56297,-0.350015), (56298,-0.107955), (56299,0.157792), (56300,-0.028416), (56301,-0.075734), (56302,-0.239181), (56303,-0.208002), (56304,-0.379808), (56305,-0.475435), (56306,-0.257997), (56307,0.054199), (56308,-0.070694), (56309,-0.103617), (56310,-0.221541), (56311,-0.053338), (56312,-0.275307), (56313,-0.295223), (56314,-0.062920), (56315,0.217229), (56316,0.061678), (56317,0.006921), (56318,-0.194609), (56319,-0.194087), (56320,-0.271599), (56321,-0.364909), (56322,-0.133995), (56323,0.137325), (56324,0.017077), (56325,-0.033033), (56326,-0.095216), (56327,0.077169), (56328,-0.250246), (56329,-0.327757), (56330,-0.072229), (56331,0.160074), (56332,0.042150), (56333,-0.001918), (56334,-0.194163), (56335,-0.191318), (56336,-0.357551), (56337,-0.385364), (56338,-0.151671), (56339,0.101071), (56340,-0.054010), (56341,-0.113876), (56342,-0.197894), (56343,-0.034794), (56344,-0.211247), (56345,-0.371907), (56346,-0.067607), (56347,0.167020), (56348,0.088581), (56349,-0.040495), (56350,-0.001421), (56351,-0.203421), (56352,-0.224264), (56353,-0.405362), (56354,-0.113598), (56355,0.159582), (56356,0.097392), (56357,-0.059085), (56358,0.114690), (56359,0.029746), (56360,-0.319034), (56361,-0.502912), (56362,0.214320), (56363,0.032295), (56364,0.000306), (56365,-0.151062), (56366,-0.186307), (56367,-0.274044), (56368,-0.400328), (56369,-0.482486), (56370,0.186444), (56371,0.006279), (56372,-0.048478), (56373,-0.174298), (56374,0.071010), (56375,-0.080821), (56376,-0.283284), (56377,-0.418860), (56378,0.230558), (56379,0.047143), (56380,0.034659), (56381,-0.116246), (56382,-0.112475), (56383,-0.298213), (56384,-0.380377), (56385,-0.519203), (56386,0.141831), (56387,0.027157), (56388,-0.008552), (56389,-0.149701), (56390,0.034294), (56391,-0.083168), (56392,-0.245218), (56393,-0.406342), (56394,0.264448), (56395,0.087069), (56396,0.023026), (56397,-0.119056), (56398,-0.125034), (56399,-0.260147), (56400,-0.315830), (56401,-0.462089), (56402,0.202195), (56403,0.050827), (56404,-0.007643), (56405,-0.156688), (56406,0.093268), (56407,-0.048814), (56408,-0.073371), (56409,-0.216843), (56410,0.044258), (56411,0.250087), (56412,0.235280), (56413,0.077406), (56414,0.065385), (56415,-0.113854), (56416,-0.107759), (56417,-0.237756), (56418,0.017772), (56419,0.244039), (56420,0.204611), (56421,0.062535), (56422,0.212623), (56423,0.119776), (56424,-0.189981), (56425,-0.339026), (56426,0.327112), (56427,0.209651), (56428,0.130279), (56429,-0.022942), (56430,-0.050755), (56431,-0.171002), (56432,-0.268958), (56433,-0.394779), (56434,0.272755), (56435,0.132075), (56436,0.049448), (56437,-0.062440), (56438,0.129457), (56439,-0.000546), (56440,-0.217875), (56441,-0.371566), (56442,0.271353), (56443,0.104656), (56444,0.067551), (56445,-0.086603), (56446,-0.068430), (56447,-0.240236), (56448,-0.549066), (56449,-0.683253), (56450,-0.024542), (56451,-0.194951), (56452,-0.223691), (56453,-0.369956), (56454,-0.141365), (56455,-0.265796), (56456,-0.420413), (56457,-0.561562), (56458,0.087393), (56459,-0.084413), (56460,-0.168894), (56461,-0.304470), (56462,-0.283974), (56463,-0.407941), (56464,-0.474307), (56465,-0.618242), (56466,0.021427), (56467,-0.135051), (56468,-0.194917), (56469,-0.304012), (56470,-0.066136), (56471,-0.227723), (56472,-0.482208), (56473,-0.511881), (56474,-0.293509), (56475,-0.046347), (56476,-0.177277), (56477,-0.238533), (56478,-0.445636), (56479,-0.441402), (56480,-0.575582), (56481,-0.625229), (56482,-0.384566), (56483,-0.093271), (56484,-0.272040), (56485,-0.277562), (56486,-0.371792), (56487,-0.208235), (56488,-0.395370), (56489,-0.477991), (56490,-0.236402), (56491,0.051180), (56492,-0.114590), (56493,-0.140079), (56494,-0.338823), (56495,-0.282567), (56496,-0.463196), (56497,-0.518416), (56498,-0.236877), (56499,0.022371), (56500,-0.106699), (56501,-0.165639), (56502,-0.227359), (56503,-0.073551), (56504,-0.444166), (56505,-0.497989), (56506,-0.255467), (56507,0.020036), (56508,-0.119253), (56509,-0.157285), (56510,-0.343493), (56511,-0.322070), (56512,-0.487834), (56513,-0.532835), (56514,-0.314000), (56515,-0.030138), (56516,-0.171750), (56517,-0.233940), (56518,-0.308201), (56519,-0.165540), (56520,-0.348498), (56521,-0.370268), (56522,-0.157940), (56523,0.133355), (56524,-0.023586), (56525,-0.066727), (56526,-0.268727), (56527,-0.265883), (56528,-0.423757), (56529,-0.473397), (56530,-0.210900), (56531,0.042768), (56532,-0.136934), (56533,-0.173576), (56534,-0.231576), (56535,-0.059660), (56536,-0.515270), (56537,-0.549589), (56538,-0.275476), (56539,-0.025991), (56540,-0.200113), (56541,-0.230719), (56542,-0.418317), (56543,-0.408503), (56544,-0.577986), (56545,-0.607195), (56546,-0.338192), (56547,-0.082664), (56548,-0.229392), (56549,-0.314336), (56550,-0.385812), (56551,-0.234791), (56552,-0.376873), (56553,-0.387961), (56554,-0.185851), (56555,0.139350), (56556,-0.027809), (56557,-0.069091), (56558,-0.288743), (56559,-0.276606), (56560,-0.460491), (56561,-0.526393), (56562,-0.281084), (56563,0.003711), (56564,-0.203862), (56565,-0.241430), (56566,-0.340776), (56567,-0.130301), (56568,-0.344380), (56569,-0.423751), (56570,-0.136633), (56571,0.140260), (56572,0.006544), (56573,-0.021269), (56574,-0.254390), (56575,-0.259904), (56576,-0.411272), (56577,-0.458596), (56578,-0.171948), (56579,0.106805), (56580,-0.030625), (56581,-0.096991), (56582,-0.202373), (56583,-0.067151), (56584,-0.398279), (56585,-0.453962), (56586,-0.238377), (56587,0.068709), (56588,-0.079409), (56589,-0.125800), (56590,-0.282741), (56591,-0.323565), (56592,-0.479110), (56593,-0.507856), (56594,-0.237926), (56595,0.035254), (56596,-0.091493), (56597,-0.178297), (56598,-0.237700), (56599,-0.105727), (56600,-0.229688), (56601,-0.372233), (56602,-0.092084), (56603,0.147188), (56604,0.129131), (56605,-0.012017), (56606,-0.030544), (56607,-0.230221), (56608,-0.281258), (56609,-0.439126), (56610,-0.158050), (56611,0.081223), (56612,0.020893), (56613,-0.144414), (56614,-0.038452), (56615,-0.135938), (56616,-0.429903), (56617,-0.565479), (56618,0.119242), (56619,-0.042808), (56620,-0.139368), (56621,-0.273084), (56622,-0.293001), (56623,-0.458771), (56624,-0.508418), (56625,-0.627269), (56626,0.056990), (56627,-0.098098), (56628,-0.150988), (56629,-0.315368), (56630,-0.071449), (56631,-0.215848), (56632,-0.374649), (56633,-0.482354), (56634,0.180997), (56635,0.017556), (56636,0.011108), (56637,-0.171850), (56638,-0.207089), (56639,-0.364036), (56640,-0.405781), (56641,-0.545077), (56642,0.108061), (56643,-0.027515), (56644,-0.120355), (56645,-0.285661), (56646,-0.009226), (56647,-0.189397), (56648,-0.353301), (56649,-0.535326), (56650,0.146139), (56651,0.018459), (56652,-0.041401), (56653,-0.195092), (56654,-0.200143), (56655,-0.358480), (56656,-0.416024), (56657,-0.596652), (56658,0.128013), (56659,-0.036824), (56660,-0.097147), (56661,-0.235980), (56662,-0.004140), (56663,-0.154575), (56664,-0.188893), (56665,-0.362559), (56666,-0.085660), (56667,0.130382), (56668,0.108612), (56669,-0.048799), (56670,-0.015760), (56671,-0.161556), (56672,-0.233031), (56673,-0.400191), (56674,-0.139553), (56675,0.076958), (56676,0.055645), (56677,-0.083644), (56678,0.076199), (56679,0.016339), (56680,-0.237219), (56681,-0.396483), (56682,0.252472), (56683,0.110853), (56684,0.040311), (56685,-0.088765), (56686,-0.123078), (56687,-0.258190), (56688,-0.305978), (56689,-0.468955), (56690,0.168385), (56691,0.036528), (56692,-0.030301), (56693,-0.153805), (56694,0.082218), (56695,-0.065437), (56696,-0.280442), (56697,-0.483369), (56698,0.187884), (56699,0.072746), (56700,-0.024740), (56701,-0.167749), (56702,-0.169550), (56703,-0.334387), (56704,-0.610244), (56705,-0.765788), (56706,-0.089426), (56707,-0.269134), (56708,-0.263503), (56709,-0.401396), (56710,-0.215542), (56711,-0.342758), (56712,-0.489017), (56713,-0.687297), (56714,0.001601), (56715,-0.159059), (56716,-0.191048), (56717,-0.301077), (56718,-0.310775), (56719,-0.480721), (56720,-0.522009), (56721,-0.660835), (56722,-0.008630), (56723,-0.163248), (56724,-0.235186), (56725,-0.401883), (56726,-0.172366), (56727,-0.317234), (56728,-0.292555), (56729,-0.383542), (56730,-0.568354), (56731,0.103363), (56732,-0.061474), (56733,-0.109725), (56734,-0.235082), (56735,-0.245713), (56736,-0.373386), (56737,-0.446722), (56738,-0.602272), (56739,0.120539), (56740,-0.068455), (56741,-0.131102), (56742,-0.315450), (56743,-0.071537), (56744,-0.483021), (56745,-0.499219), (56746,-0.261806), (56747,0.030416), (56748,-0.127922), (56749,-0.232371), (56750,-0.392104), (56751,-0.398083), (56752,-0.564779), (56753,-0.600958), (56754,-0.350069), (56755,-0.054598), (56756,-0.202710), (56757,-0.270936), (56758,-0.349844), (56759,-0.250388), (56760,-0.544353), (56761,-0.587958), (56762,-0.368196), (56763,-0.094090), (56764,-0.217587), (56765,-0.267228), (56766,-0.423705), (56767,-0.423184), (56768,-0.553651), (56769,-0.645101), (56770,-0.415584), (56771,-0.121039), (56772,-0.283553), (56773,-0.343883), (56774,-0.378665), (56775,-0.247619), (56776,-0.493745), (56777,-0.525740), (56778,-0.243268), (56779,0.059172), (56780,-0.143754), (56781,-0.224052), (56782,-0.387036), (56783,-0.352607), (56784,-0.498396), (56785,-0.566158), (56786,-0.316667), (56787,-0.061139), (56788,-0.220866), (56789,-0.264477), (56790,-0.354067), (56791,-0.216052), (56792,-0.385535), (56793,-0.424030), (56794,-0.569825), (56795,0.083306), (56796,-0.109401), (56797,-0.163688), (56798,-0.320629), (56799,-0.306639), (56800,-0.445001), (56801,-0.502544), (56802,-0.630688), (56803,0.061466), (56804,-0.073646), (56805,-0.168809), (56806,-0.326677), (56807,-0.076259), (56808,-0.237382), (56809,-0.306071), (56810,-0.468585), (56811,0.218923), (56812,0.066159), (56813,-0.006713), (56814,-0.165513), (56815,-0.171028), (56816,-0.334475), (56817,-0.388299), (56818,-0.565678), (56819,0.119971), (56820,-0.031397), (56821,-0.065709), (56822,-0.213364), (56823,0.011976), (56824,-0.143111), (56825,-0.200185), (56826,-0.371991), (56827,0.316907), (56828,0.146498), (56829,0.060621), (56830,-0.071236), (56831,-0.050277), (56832,-0.196535), (56833,-0.271730), (56834,-0.471870), (56835,0.205882), (56836,0.082385), (56837,0.017879), (56838,-0.133026), (56839,0.094632), (56840,-0.215125), (56841,-0.264309), (56842,-0.429146), (56843,0.272295), (56844,0.105598), (56845,0.045738), (56846,-0.139074), (56847,-0.142735), (56848,-0.267629), (56849,-0.346067), (56850,-0.486753), (56851,0.178458), (56852,0.023377), (56853,-0.008619), (56854,-0.140945), (56855,0.099724), (56856,-0.289005), (56857,-0.445019), (56858,-0.147682), (56859,0.067433), (56860,-0.004969), (56861,-0.176775), (56862,-0.144670), (56863,-0.305794), (56864,-0.345679), (56865,-0.491474), (56866,-0.219227), (56867,0.039093), (56868,-0.030065), (56869,-0.144733), (56870,0.018360), (56871,-0.073554), (56872,-0.166394), (56873,-0.333090), (56874,-0.050625), (56875,0.164960), (56876,0.152006), (56877,-0.056957), (56878,-0.001163), (56879,-0.203620), (56880,-0.248158), (56881,-0.388380), (56882,-0.106835), (56883,0.141260), (56884,0.082327), (56885,-0.082516), (56886,0.071291), (56887,0.005852), (56888,-0.152949), (56889,-0.259258), (56890,-0.036246), (56891,0.187698), (56892,0.151062), (56893,-0.020744), (56894,-0.046240), (56895,-0.188315), (56896,-0.252358), (56897,-0.432060), (56898,-0.125437), (56899,0.113366), (56900,0.060476), (56901,-0.075101), (56902,0.047580), (56903,-0.031792), (56904,-0.165971), (56905,-0.334528), (56906,-0.072494), (56907,0.179785), (56908,0.138033), (56909,0.019182), (56910,-0.039751), (56911,-0.180906), (56912,-0.219865), (56913,-0.381452), (56914,-0.103163), (56915,0.115209), (56916,0.056739), (56917,-0.110421), (56918,0.069854), (56919,-0.050393), (56920,-0.284904), (56921,-0.447418), (56922,-0.174238), (56923,0.039950), (56924,-0.020379), (56925,-0.158742), (56926,-0.117344), (56927,-0.263139), (56928,-0.355979), (56929,-0.527322), (56930,-0.229528), (56931,0.004172), (56932,-0.058944), (56933,-0.191264), (56934,-0.057901), (56935,-0.120084), (56936,-0.404300), (56937,-0.557528), (56938,0.154601), (56939,0.008343), (56940,-0.009251), (56941,-0.199172), (56942,-0.230704), (56943,-0.375566), (56944,-0.457260), (56945,-0.591446), (56946,0.106751), (56947,-0.029289), (56948,-0.062211), (56949,-0.181532), (56950,0.011292), (56951,-0.124748), (56952,-0.362514), (56953,-0.506913), (56954,0.117421), (56955,-0.029764), (56956,-0.095666), (56957,-0.200585), (56958,-0.214929), (56959,-0.358865), (56960,-0.392720), (56961,-0.460476), (56962,-0.228636), (56963,0.062196), (56964,-0.145377), (56965,-0.202457), (56966,-0.272536), (56967,-0.092254), (56968,-0.336521), (56969,-0.387094), (56970,-0.191021), (56971,0.118389), (56972,-0.095690), (56973,-0.076584), (56974,-0.303205), (56975,-0.298037), (56976,-0.474026), (56977,-0.512521), (56978,-0.254207), (56979,0.017583), (56980,-0.154687), (56981,-0.169494), (56982,-0.233073), (56983,-0.084382), (56984,-0.452203), (56985,-0.528325), (56986,-0.316460), (56987,-0.039097), (56988,-0.208580), (56989,-0.279129), (56990,-0.417955), (56991,-0.394672), (56992,-0.532571), (56993,-0.578036), (56994,-0.330404), (56995,-0.092521), (56996,-0.261541), (56997,-0.270312), (56998,-0.324599), (56999,-0.202382), (57000,-0.281290), (57001,-0.407110), (57002,-0.064257), (57003,-0.261147), (57004,-0.012582), (57005,-0.146768), (57006,-0.221956), (57007,-0.358459), (57008,-0.344006), (57009,-0.500947), (57010,-0.163203), (57011,-0.305285), (57012,0.006448), (57013,-0.156529), (57014,-0.130930), (57015,-0.292980), (57016,-0.265978), (57017,-0.412243), (57018,-0.085645), (57019,-0.256055), (57020,0.019911), (57021,-0.147718), (57022,-0.244741), (57023,-0.421187), (57024,-0.371894), (57025,-0.546956), (57026,-0.151611), (57027,-0.312271), (57028,-0.050237), (57029,-0.220653), (57030,-0.193651), (57031,-0.374750), (57032,-0.223266), (57033,-0.356519), (57034,-0.031781), (57035,-0.239817), (57036,0.056118), (57037,-0.111969), (57038,-0.211315), (57039,-0.334812), (57040,-0.326395), (57041,-0.485195), (57042,-0.137696), (57043,-0.288601), (57044,0.039387), (57045,-0.127309), (57046,-0.093344), (57047,-0.248895), (57048,-0.358923), (57049,-0.488457), (57050,-0.191589), (57051,-0.352250), (57052,-0.085570), (57053,-0.206281), (57054,-0.297267), (57055,-0.457928), (57056,-0.468089), (57057,-0.653364), (57058,-0.288676), (57059,-0.414033), (57060,-0.106483), (57061,-0.269930), (57062,-0.220173), (57063,-0.396155), (57064,-0.264183), (57065,-0.412301), (57066,-0.097782), (57067,-0.265875), (57068,0.030999), (57069,-0.124552), (57070,-0.194167), (57071,-0.337176), (57072,-0.356166), (57073,-0.501028), (57074,-0.147956), (57075,-0.292824), (57076,0.017982), (57077,-0.140355), (57078,-0.109640), (57079,-0.267514), (57080,-0.194996), (57081,-0.336608), (57082,0.017860), (57083,-0.151159), (57084,0.184261), (57085,0.047289), (57086,-0.036729), (57087,-0.161616), (57088,-0.231701), (57089,-0.403044), (57090,-0.036496), (57091,-0.191584), (57092,0.069987), (57093,-0.076742), (57094,-0.025588), (57095,-0.182066), (57096,-0.187117), (57097,-0.351961), (57098,-0.022106), (57099,-0.175797), (57100,0.089017), (57101,-0.057242), (57102,-0.123608), (57103,-0.307493), (57104,-0.276314), (57105,-0.396562), (57106,-0.066714), (57107,-0.210186), (57108,0.082969), (57109,-0.055857), (57110,-0.009814), (57111,-0.183479), (57112,-0.145801), (57113,-0.230745), (57114,-0.349133), (57115,0.346734), (57116,0.147991), (57117,0.071406), (57118,-0.089255), (57119,-0.062722), (57120,-0.212231), (57121,-0.300894), (57122,-0.422068), (57123,0.228746), (57124,0.069013), (57125,0.023548), (57126,-0.167299), (57127,0.045962), (57128,-0.309323), (57129,-0.406346), (57130,-0.143386), (57131,0.139550), (57132,-0.004849), (57133,-0.018730), (57134,-0.212827), (57135,-0.187691), (57136,-0.337663), (57137,-0.387310), (57138,-0.135495), (57139,0.114923), (57140,-0.032732), (57141,-0.062398), (57142,-0.155708), (57143,-0.019552), (57144,-0.281470), (57145,-0.296740), (57146,-0.100667), (57147,0.169257), (57148,0.041576), (57149,0.008654), (57150,-0.182194), (57151,-0.215579), (57152,-0.386922), (57153,-0.412412), (57154,-0.160133), (57155,0.134411), (57156,0.024383), (57157,-0.029441), (57158,-0.090234), (57159,0.024550), (57160,-0.198814), (57161,-0.266570), (57162,-0.038913), (57163,0.228694), (57164,0.066180), (57165,0.006777), (57166,-0.178034), (57167,-0.119912), (57168,-0.289401), (57169,-0.378992), (57170,-0.138786), (57171,0.166904), (57172,-0.006292), (57173,-0.074981), (57174,-0.132524), (57175,0.016637), (57176,-0.139840), (57177,-0.230364), (57178,-0.343179), (57179,0.315069), (57180,0.209223), (57181,0.172118), (57182,-0.029882), (57183,-0.067450), (57184,-0.151461), (57185,-0.212254), (57186,-0.385920), (57187,0.281150), (57188,0.117703), (57189,0.087104), (57190,-0.095384), (57191,0.147602), (57192,-0.224403), (57193,-0.277763), (57194,-0.021765), (57195,0.307619), (57196,0.136740), (57197,0.055509), (57198,-0.147881), (57199,-0.123672), (57200,-0.292692), (57201,-0.338619), (57202,-0.087738), (57203,0.230501), (57204,0.042903), (57205,-0.000238), (57206,-0.092615), (57207,0.072338), (57208,-0.285734), (57209,-0.327016), (57210,-0.075671), (57211,0.210984), (57212,0.048464), (57213,0.014152), (57214,-0.185988), (57215,-0.204052), (57216,-0.226755), (57217,0.126787), (57218,-0.039446), (57219,0.233270), (57220,0.071214), (57221,0.086600), (57222,-0.074060), (57223,0.073711), (57224,-0.058152), (57225,0.270769), (57226,0.118004), (57227,0.367033), (57228,0.252822), (57229,0.191102), (57230,0.010473), (57231,0.028640), (57232,-0.123191), (57233,0.200620), (57234,0.075726), (57235,0.325218), (57236,0.190105), (57237,0.200383), (57238,0.034149), (57239,0.211181), (57240,-0.043311), (57241,0.225229), (57242,0.188588), (57243,0.006099), (57244,0.324331), (57245,0.148812), (57246,0.096379), (57247,-0.094006), (57248,-0.069327), (57249,0.185738), (57250,0.117512), (57251,-0.059403), (57252,0.262085), (57253,0.204078), (57254,0.166510), (57255,-0.027594), (57256,0.077441), (57257,0.306958), (57258,0.252671), (57259,0.119418), (57260,0.367050), (57261,0.191061), (57262,0.158139), (57263,0.026276), (57264,0.010079), (57265,0.240059), (57266,0.168584), (57267,0.021862), (57268,0.322912), (57269,0.248181), (57270,0.210619), (57271,0.008619), (57272,-0.091190), (57273,0.180593), (57274,0.152317), (57275,0.003735), (57276,0.242545), (57277,0.072592), (57278,0.055468), (57279,-0.127027), (57280,-0.109781), (57281,0.079324), (57282,0.049188), (57283,-0.119362), (57284,0.164963), (57285,0.070727), (57286,0.020616), (57287,-0.107527), (57288,0.126173), (57289,0.334788), (57290,0.289324), (57291,0.159321), (57292,0.446902), (57293,0.247689), (57294,0.217089), (57295,0.056429), (57296,0.084821), (57297,0.348245), (57298,0.302781), (57299,0.115646), (57300,0.429702), (57301,0.339648), (57302,0.285361), (57303,0.127951), (57304,0.040220), (57305,0.242799), (57306,0.252607), (57307,0.084984), (57308,0.389284), (57309,0.217014), (57310,0.153898), (57311,-0.031377), (57312,-0.013210), (57313,0.210734), (57314,0.158307), (57315,-0.010713), (57316,0.265717), (57317,0.190058), (57318,0.105114), (57319,-0.047644), (57320,0.096401), (57321,0.313846), (57322,0.224719), (57323,0.107258), (57324,0.379511), (57325,0.196553), (57326,0.135760), (57327,-0.059734), (57328,-0.025769), (57329,0.229295), (57330,0.189404), (57331,0.047791), (57332,0.367420), (57333,0.292232), (57334,0.246304), (57335,0.046627), (57336,0.308191), (57337,0.156823), (57338,0.454161), (57339,0.335767), (57340,0.663761), (57341,0.505424), (57342,0.429765), (57343,0.258423), (57344,0.280779), (57345,0.153562), (57346,0.466221), (57347,0.288842), (57348,0.587106), (57349,0.447354), (57350,0.469703), (57351,0.300220), (57352,0.259865), (57353,0.122893), (57354,0.464356), (57355,0.264679), (57356,0.585241), (57357,0.446409), (57358,0.328484), (57359,0.230071), (57360,0.234306), (57361,0.086188), (57362,0.429511), (57363,0.291148), (57364,0.549926), (57365,0.413423), (57366,0.410225), (57367,0.271399), (57368,0.197601), (57369,0.180471), (57370,0.426249), (57371,0.690136), (57372,0.546664), (57373,0.515139), (57374,0.353082), (57375,0.351286), (57376,0.158109), (57377,0.093603), (57378,0.327766), (57379,0.611628), (57380,0.460260), (57381,0.455209), (57382,0.377691), (57383,0.485976), (57384,0.034542), (57385,0.386224), (57386,0.222778), (57387,0.462050), (57388,0.356205), (57389,0.296802), (57390,0.100844), (57391,0.086501), (57392,0.000623), (57393,0.309570), (57394,0.180500), (57395,0.427668), (57396,0.258649), (57397,0.271712), (57398,0.130100), (57399,0.276931), (57400,0.143678), (57401,0.085208), (57402,0.337023), (57403,0.609740), (57404,0.478346), (57405,0.435205), (57406,0.236918), (57407,0.282499), (57408,0.124161), (57409,0.054083), (57410,0.318897), (57411,0.545627), (57412,0.429562), (57413,0.411036), (57414,0.294044), (57415,0.484075), (57416,0.180818), (57417,0.167870), (57418,0.441513), (57419,0.684499), (57420,0.538710), (57421,0.444474), (57422,0.255479), (57423,0.305700), (57424,0.112065), (57425,0.068924), (57426,0.298905), (57427,0.587413), (57428,0.439295), (57429,0.414268), (57430,0.353012), (57431,0.510532), (57432,0.196593), (57433,0.171103), (57434,0.411302), (57435,0.653825), (57436,0.511749), (57437,0.489509), (57438,0.314917), (57439,0.333553), (57440,0.177539), (57441,0.107923), (57442,0.313746), (57443,0.601791), (57444,0.460642), (57445,0.400782), (57446,0.323728), (57447,0.461743), (57448,0.129218), (57449,0.444207), (57450,0.318850), (57451,0.597603), (57452,0.465740), (57453,0.351535), (57454,0.170437), (57455,0.170495), (57456,0.012621), (57457,0.376375), (57458,0.216185), (57459,0.489364), (57460,0.364934), (57461,0.394259), (57462,0.264719), (57463,0.416203), (57464,0.013079), (57465,0.358255), (57466,0.211527), (57467,0.499572), (57468,0.295255), (57469,0.229353), (57470,0.079375), (57471,0.127741), (57472,-0.077045), (57473,0.178946), (57474,0.303486), (57475,0.140509), (57476,0.091795), (57477,0.033789), (57478,0.301395), (57479,0.158387), (57480,0.000049), (57481,0.351732), (57482,0.186889), (57483,0.157223), (57484,0.030932), (57485,-0.081419), (57486,-0.248579), (57487,0.043649), (57488,-0.123518), (57489,0.249066), (57490,0.115813), (57491,0.279839), (57492,0.103387), (57493,0.120164), (57494,0.007349), (57495,0.255444), (57496,0.068773), (57497,0.063258), (57498,0.296488), (57499,0.251030), (57500,0.080614), (57501,0.035150), (57502,-0.092061), (57503,0.225708), (57504,0.046933), (57505,0.002402), (57506,0.262576), (57507,0.388969), (57508,0.206017), (57509,0.168912), (57510,0.081645), (57511,0.337643), (57512,0.020447), (57513,0.344722), (57514,0.216115), (57515,0.231502), (57516,0.085706), (57517,-0.001567), (57518,-0.135747), (57519,0.149048), (57520,-0.018118), (57521,0.341924), (57522,0.137137), (57523,0.267720), (57524,0.095450), (57525,0.151243), (57526,0.017990), (57527,0.264696), (57528,-0.146788), (57529,0.220680), (57530,0.110188), (57531,0.136720), (57532,-0.055061), (57533,-0.086587), (57534,-0.226346), (57535,0.025933), (57536,-0.109174), (57537,0.198376), (57538,0.094384), (57539,0.228216), (57540,0.056410), (57541,0.102917), (57542,-0.038695), (57543,0.226589), (57544,0.036661), (57545,0.381374), (57546,0.206782), (57547,0.153421), (57548,-0.003056), (57549,-0.072672), (57550,-0.178054), (57551,0.090480), (57552,-0.039987), (57553,0.318195), (57554,0.136170), (57555,0.292763), (57556,0.140926), (57557,0.162818), (57558,-0.020140), (57559,0.296702), (57560,0.124896), (57561,0.016727), (57562,0.284798), (57563,0.285782), (57564,0.123269), (57565,0.096383), (57566,-0.098185), (57567,0.149447), (57568,0.036169), (57569,0.019039), (57570,0.258311), (57571,0.317824), (57572,0.216155), (57573,0.156295), (57574,0.101075), (57575,0.396552), (57576,0.235429), (57577,0.204360), (57578,0.424591), (57579,0.414893), (57580,0.283963), (57581,0.219451), (57582,0.053687), (57583,0.342659), (57584,0.144842), (57585,0.097054), (57586,0.324248), (57587,0.479909), (57588,0.375923), (57589,0.337428), (57590,0.209284), (57591,0.514511), (57592,0.256307), (57593,0.216885), (57594,0.447329), (57595,0.486403), (57596,0.315530), (57597,0.254737), (57598,0.069925), (57599,0.343568), (57600,0.215425), (57601,0.133267), (57602,0.405051), (57603,0.567680), (57604,0.435354), (57605,0.391286), (57606,0.307269), (57607,0.613892), (57608,0.265582), (57609,0.207575), (57610,0.412008), (57611,0.456655), (57612,0.302038), (57613,0.269579), (57614,0.040178), (57615,0.344941), (57616,0.237236), (57617,0.192235), (57618,0.430111), (57619,0.549548), (57620,0.412112), (57621,0.338314), (57622,0.301679), (57623,0.591113), (57624,0.179160), (57625,0.064028), (57626,0.448684), (57627,0.309389), (57628,0.219798), (57629,0.049389), (57630,0.264040), (57631,0.121501), (57632,0.068604), (57633,-0.115281), (57634,0.461678), (57635,0.321925), (57636,0.281570), (57637,0.102795), (57638,0.478629), (57639,0.346302), (57640,0.260431), (57641,0.097911), (57642,0.488610), (57643,0.365576), (57644,0.318252), (57645,0.185932), (57646,0.394078), (57647,0.203230), (57648,0.171235), (57649,0.052384), (57650,0.568491), (57651,0.411550), (57652,0.364696), (57653,0.225400), (57654,0.576613), (57655,0.432214), (57656,0.274346), (57657,0.117399), (57658,0.537359), (57659,0.394356), (57660,0.347496), (57661,0.147819), (57662,0.367117), (57663,0.235260), (57664,0.155426), (57665,0.007771), (57666,0.569401), (57667,0.408740), (57668,0.368855), (57669,0.243035), (57670,0.577522), (57671,0.399217), (57672,0.250172), (57673,0.128528), (57674,0.513654), (57675,0.338591), (57676,0.296383), (57677,0.196110), (57678,0.409829), (57679,0.249175), (57680,0.206034), (57681,0.028655), (57682,0.568914), (57683,0.394791), (57684,0.345607), (57685,0.232329), (57686,0.591901), (57687,0.460971), (57688,0.192553), (57689,0.023534), (57690,0.415159), (57691,0.280979), (57692,0.202998), (57693,0.080428), (57694,0.316450), (57695,0.161363), (57696,0.123795), (57697,0.007730), (57698,0.496900), (57699,0.345995), (57700,0.325615), (57701,0.184003), (57702,0.529179), (57703,0.376878), (57704,0.217151), (57705,0.541889), (57706,0.400277), (57707,0.427736), (57708,0.253606), (57709,0.175162), (57710,0.033086), (57711,0.332740), (57712,0.197634), (57713,0.515403), (57714,0.335701), (57715,0.498794), (57716,0.391089), (57717,0.385104), (57718,0.218877), (57719,0.462790), (57720,0.077316), (57721,0.342600), (57722,0.343122), (57723,0.199650), (57724,0.126778), (57725,-0.047815), (57726,0.219792), (57727,0.052169), (57728,0.010418), (57729,-0.036437), (57730,0.192617), (57731,0.344095), (57732,0.196446), (57733,0.158414), (57734,0.065568), (57735,0.351290), (57736,-0.008636), (57737,0.335614), (57738,0.197251), (57739,0.195449), (57740,0.039435), (57741,-0.010675), (57742,-0.153684), (57743,0.152939), (57744,-0.047664), (57745,0.260355), (57746,0.147541), (57747,0.283226), (57748,0.124426), (57749,0.128667), (57750,-0.003660), (57751,0.265337), (57752,0.227305), (57753,0.104741), (57754,0.478252), (57755,0.303189), (57756,0.287919), (57757,0.147697), (57758,0.078544), (57759,-0.054709), (57760,0.207325), (57761,0.019727), (57762,0.350038), (57763,0.178696), (57764,0.341789), (57765,0.163020), (57766,0.223922), (57767,0.079987), (57768,0.067039), (57769,0.326281), (57770,0.300791), (57771,0.135491), (57772,0.172706), (57773,-0.019075), (57774,-0.078472), (57775,-0.221017), (57776,0.037297), (57777,0.275180), (57778,0.224143), (57779,0.095993), (57780,0.269775), (57781,0.191794), (57782,0.136580), (57783,0.000534), (57784,0.217515), (57785,0.108877), (57786,0.417360), (57787,0.252053), (57788,0.271159), (57789,0.082165), (57790,0.015336), (57791,-0.175055), (57792,0.118563), (57793,-0.046274), (57794,0.303548), (57795,0.144748), (57796,0.283226), (57797,0.153687), (57798,0.143526), (57799,0.017242), (57800,0.125057), (57801,0.361543), (57802,0.354169), (57803,0.185149), (57804,0.203785), (57805,0.002718), (57806,-0.021381), (57807,-0.187614), (57808,0.115296), (57809,0.357818), (57810,0.266831), (57811,0.098275), (57812,0.266484), (57813,0.204295), (57814,0.140252), (57815,0.012572), (57816,0.270423), (57817,0.090721), (57818,0.420569), (57819,0.278957), (57820,0.331963), (57821,0.142042), (57822,0.028301), (57823,-0.130500), (57824,0.114809), (57825,-0.014261), (57826,0.348560), (57827,0.204162), (57828,0.354713), (57829,0.184766), (57830,0.221054), (57831,0.070150), (57832,0.352158), (57833,0.172450), (57834,0.487902), (57835,0.336534), (57836,0.318007), (57837,0.199620), (57838,0.132327), (57839,-0.014395), (57840,0.266211), (57841,0.120886), (57842,0.430296), (57843,0.313761), (57844,0.468958), (57845,0.286007), (57846,0.352488), (57847,0.191828), (57848,0.398121), (57849,0.236533), (57850,0.557089), (57851,0.431732), (57852,0.453624), (57853,0.275776), (57854,0.195478), (57855,0.029244), (57856,0.303351), (57857,0.180780), (57858,0.538499), (57859,0.413142), (57860,0.557193), (57861,0.374705), (57862,0.413779), (57863,0.218749), (57864,0.317278), (57865,0.222114), (57866,0.566827), (57867,0.439147), (57868,0.454997), (57869,0.288301), (57870,0.207996), (57871,0.051519), (57872,0.340490), (57873,0.181690), (57874,0.518970), (57875,0.366212), (57876,0.513050), (57877,0.360286), (57878,0.407256), (57879,0.263784), (57880,0.245727), (57881,0.160313), (57882,0.441858), (57883,0.436801), (57884,0.236197), (57885,0.190269), (57886,-0.000115), (57887,0.273065), (57888,0.111014), (57889,0.040002), (57890,0.295994), (57891,0.500896), (57892,0.333730), (57893,0.263187), (57894,0.194035), (57895,0.511804), (57896,0.293549), (57897,0.242975), (57898,0.452517), (57899,0.493915), (57900,0.317463), (57901,0.271535), (57902,0.115521), (57903,0.383591), (57904,0.241515), (57905,0.166320), (57906,0.429281), (57907,0.544072), (57908,0.395490), (57909,0.367677), (57910,0.296665), (57911,0.555913), (57912,0.284703), (57913,0.248061), (57914,0.470152), (57915,0.515726), (57916,0.315122), (57917,0.265475), (57918,0.083920), (57919,0.315290), (57920,0.168568), (57921,0.136573), (57922,0.389784), (57923,0.563560), (57924,0.395003), (57925,0.336997), (57926,0.254376), (57927,0.505257), (57928,0.293045), (57929,0.215527), (57930,0.412997), (57931,0.479009), (57932,0.350402), (57933,0.301225), (57934,0.160076), (57935,0.441615), (57936,0.258193), (57937,0.200193), (57938,0.435746), (57939,0.609058), (57940,0.427033), (57941,0.374606), (57942,0.287332), (57943,0.564695), (57944,0.221025), (57945,0.158378), (57946,0.401364), (57947,0.410708), (57948,0.255164), (57949,0.211553), (57950,0.045789), (57951,0.312926), (57952,0.190825), (57953,0.120740), (57954,0.363732), (57955,0.518460), (57956,0.355019), (57957,0.311878), (57958,0.218568), (57959,0.461554), (57960,0.073764), (57961,0.452378), (57962,0.298223), (57963,0.343804), (57964,0.175711), (57965,0.094016), (57966,-0.046200), (57967,0.228833), (57968,0.089081), (57969,0.405460), (57970,0.260128), (57971,0.419971), (57972,0.298791), (57973,0.275624), (57974,0.146091), (57975,0.462463), (57976,0.271616), (57977,0.176916), (57978,0.401787), (57979,0.436678), (57980,0.255586), (57981,0.215231), (57982,0.023450), (57983,0.304063), (57984,0.027743), (57985,-0.017715), (57986,0.199723), (57987,0.366066), (57988,0.212838), (57989,0.151582), (57990,0.098692), (57991,0.391840), (57992,0.183340), (57993,0.077958), (57994,0.405946), (57995,0.272693), (57996,0.272751), (57997,0.143681), (57998,0.089387), (57999,-0.102857), (58000,0.177755), (58001,0.042649), (58002,0.356235), (58003,0.216483), (58004,0.341486), (58005,0.227745), (58006,0.236162), (58007,0.033699), (58008,0.220480), (58009,0.068648), (58010,0.438439), (58011,0.254561), (58012,0.230924), (58013,0.069801), (58014,0.044781), (58015,-0.096374), (58016,0.174019), (58017,0.000823), (58018,0.349249), (58019,0.160718), (58020,0.301519), (58021,0.152474), (58022,0.222669), (58023,0.062942), (58024,0.049525), (58025,0.319918), (58026,0.267021), (58027,0.102184), (58028,0.113852), (58029,-0.064918), (58030,-0.115491), (58031,-0.269183), (58032,0.025825), (58033,0.253019), (58034,0.217774), (58035,0.085454), (58036,0.230895), (58037,0.106935), (58038,0.089805), (58039,-0.046698), (58040,0.184209), (58041,0.029591), (58042,0.381267), (58043,0.214107), (58044,0.220201), (58045,0.091594), (58046,0.001541), (58047,-0.118243), (58048,0.134962), (58049,-0.029875), (58050,0.299509), (58051,0.153251), (58052,0.283827), (58053,0.145928), (58054,0.143663), (58055,-0.037429), (58056,0.244573), (58057,0.111320), (58058,0.449990), (58059,0.291659), (58060,0.261524), (58061,0.122228), (58062,0.001054), (58063,-0.158210), (58064,0.153059), (58065,0.010977), (58066,0.273938), (58067,0.137899), (58068,0.311680), (58069,0.193286), (58070,0.228184), (58071,0.066597), (58072,0.147011), (58073,-0.009936), (58074,0.310626), (58075,0.170867), (58076,0.200655), (58077,0.046031), (58078,-0.045882), (58079,-0.180062), (58080,0.125635), (58081,-0.033166), (58082,0.351027), (58083,0.204768), (58084,0.362752), (58085,0.194659), (58086,0.214229), (58087,0.030344), (58088,0.271476), (58089,0.135430), (58090,0.498722), (58091,0.370115), (58092,0.371569), (58093,0.218342), (58094,0.131074), (58095,-0.027726), (58096,0.238484), (58097,0.102908), (58098,0.410458), (58099,0.247944), (58100,0.418470), (58101,0.278248), (58102,0.302463), (58103,0.171064), (58104,0.313255), (58105,0.133553), (58106,0.442036), (58107,0.349660), (58108,0.374332), (58109,0.225751), (58110,0.144520), (58111,-0.043078), (58112,0.205487), (58113,0.087562), (58114,0.446207), (58115,0.279511), (58116,0.428672), (58117,0.282877), (58118,0.311269), (58119,0.158504), (58120,0.304879), (58121,0.112635), (58122,0.481962), (58123,0.361715), (58124,0.315324), (58125,0.180674), (58126,0.062750), (58127,-0.077003), (58128,0.170629), (58129,0.035053), (58130,0.415996), (58131,0.243257), (58132,0.410997), (58133,0.236404), (58134,0.247608), (58135,0.127360), (58136,0.329476), (58137,0.253355), (58138,0.084799), (58139,0.481533), (58140,0.348280), (58141,0.280988), (58142,0.076202), (58143,0.373533), (58144,0.251432), (58145,0.173450), (58146,0.009540), (58147,0.553055), (58148,0.424448), (58149,0.339041), (58150,0.191849), (58151,0.571866), (58152,0.244914), (58153,0.161366), (58154,0.429436), (58155,0.402550), (58156,0.259078), (58157,0.185743), (58158,0.034839), (58159,0.285727), (58160,0.181271), (58161,0.124191), (58162,0.382512), (58163,0.509375), (58164,0.374726), (58165,0.290708), (58166,0.253140), (58167,0.530039), (58168,0.193338), (58169,0.110711), (58170,0.344874), (58171,0.347255), (58172,0.134109), (58173,0.146709), (58174,-0.050181), (58175,0.246223), (58176,0.079063), (58177,0.034989), (58178,0.274725), (58179,0.433178), (58180,0.266482), (58181,0.245632), (58182,0.118422), (58183,0.454769), (58184,0.198887), (58185,0.128808), (58186,0.349966), (58187,0.339335), (58188,0.205156), (58189,0.193598), (58190,0.011573), (58191,0.281966), (58192,0.106911), (58193,0.070275), (58194,0.275171), (58195,0.409004), (58196,0.298975), (58197,0.227500), (58198,0.123044), (58199,0.411553), (58200,0.305707), (58201,0.231439), (58202,0.078681), (58203,0.487025), (58204,0.374210), (58205,0.314350), (58206,0.117923), (58207,0.370665), (58208,0.251350), (58209,0.227251), (58210,0.050335), (58211,0.569699), (58212,0.403929), (58213,0.373793), (58214,0.237753), (58215,0.584790), (58216,0.200243), (58217,0.459491), (58218,0.412166), (58219,0.299815), (58220,0.330530), (58221,0.131317), (58222,0.108150), (58223,-0.071089), (58224,0.153782), (58225,0.429285), (58226,0.398686), (58227,0.225953), (58228,0.375577), (58229,0.318034), (58230,0.276753), (58231,0.088685), (58232,0.248065), (58233,0.161724), (58234,0.397284), (58235,0.421030), (58236,0.251547), (58237,0.227447), (58238,0.048672), (58239,0.366447), (58240,0.041355), (58241,-0.134164), (58242,0.211939), (58243,0.077760), (58244,0.233420), (58245,0.106667), (58246,0.116944), (58247,-0.046033), (58248,0.191843), (58249,0.005635), (58250,0.324337), (58251,0.192944), (58252,0.177667), (58253,0.014690), (58254,-0.033098), (58255,-0.201184), (58256,0.081745), (58257,-0.075660), (58258,0.263481), (58259,0.123722), (58260,0.274736), (58261,0.112222), (58262,0.085336), (58263,-0.031192), (58264,0.135151), (58265,-0.029222), (58266,0.270901), (58267,0.164123), (58268,0.195301), (58269,0.021635), (58270,-0.062845), (58271,-0.227219), (58272,0.079868), (58273,-0.085902), (58274,0.251848), (58275,0.090255), (58276,0.255677), (58277,0.159118), (58278,0.116440), (58279,-0.052117), (58280,0.222923), (58281,0.032538), (58282,0.412548), (58283,0.276972), (58284,0.265884), (58285,0.117766), (58286,0.039322), (58287,-0.129228), (58288,0.191327), (58289,0.065970), (58290,0.396745), (58291,0.204037), (58292,0.386642), (58293,0.242243), (58294,0.251123), (58295,0.073744), (58296,0.027347), (58297,-0.106369), (58298,0.261568), (58299,0.128315), (58300,0.113971), (58301,-0.029501), (58302,-0.120944), (58303,-0.225870), (58304,0.064498), (58305,-0.119387), (58306,0.206748), (58307,0.060953), (58308,0.211041), (58309,0.034125), (58310,0.116862), (58311,-0.039152), (58312,0.195475), (58313,0.051076), (58314,0.360022), (58315,0.224446), (58316,0.259338), (58317,0.061984), (58318,0.016520), (58319,-0.153890), (58320,0.097925), (58321,-0.013037), (58322,0.259216), (58323,0.184954), (58324,0.330396), (58325,0.177638), (58326,0.204170), (58327,-0.029883), (58328,0.097450), (58329,-0.064601), (58330,0.301007), (58331,0.152426), (58332,0.154344), (58333,-0.023499), (58334,-0.070823), (58335,-0.236123), (58336,0.037057), (58337,-0.145902), (58338,0.217390), (58339,0.083673), (58340,0.236548), (58341,0.081466), (58342,0.126114), (58343,-0.024328), (58344,-0.125997), (58345,0.179700), (58346,0.400858), (58347,0.373045), (58348,0.193343), (58349,0.204547), (58350,0.034131), (58351,0.018860), (58352,-0.178030), (58353,0.109088), (58354,0.319557), (58355,0.281062), (58356,0.126907), (58357,0.270495), (58358,0.172539), (58359,0.167024), (58360,0.427199), (58361,0.273044), (58362,0.243372), (58363,0.481718), (58364,0.448326), (58365,0.347126), (58366,0.257999), (58367,0.052286), (58368,0.386311), (58369,0.225193), (58370,0.161144), (58371,0.380442), (58372,0.550505), (58373,0.387991), (58374,0.324875), (58375,0.265942), (58376,0.056979), (58377,0.279063), (58378,0.127226), (58379,0.498883), (58380,0.349838), (58381,0.354999), (58382,0.220356), (58383,0.144234), (58384,-0.005274), (58385,0.273015), (58386,0.140226), (58387,0.466354), (58388,0.316846), (58389,0.425130), (58390,0.264007), (58391,0.291935), (58392,0.238575), (58393,0.206580), (58394,0.070077), (58395,0.451020), (58396,0.315444), (58397,0.243968), (58398,0.098173), (58399,0.349518), (58400,0.164707), (58401,0.141077), (58402,0.005501), (58403,0.520218), (58404,0.344693), (58405,0.300625), (58406,0.211034), (58407,0.554814), (58408,0.203255), (58409,0.043521), (58410,0.419354), (58411,0.283778), (58412,0.247606), (58413,0.128286), (58414,0.031732), (58415,-0.110813), (58416,0.158647), (58417,-0.008050), (58418,0.349669), (58419,0.178796), (58420,0.306586), (58421,0.099946), (58422,0.189646), (58423,0.044784), (58424,0.254326), (58425,0.194930), (58426,0.061207), (58427,0.467698), (58428,0.328408), (58429,0.295486), (58430,0.171519), (58431,0.400573), (58432,0.257101), (58433,0.151255), (58434,0.004533), (58435,0.547585), (58436,0.354408), (58437,0.340997), (58438,0.182196), (58439,0.558956), (58440,0.373218), (58441,0.219527), (58442,0.154088), (58443,0.414262), (58444,0.424076), (58445,0.254587), (58446,0.193800), (58447,0.045218), (58448,0.330470), (58449,0.168420), (58450,0.119706), (58451,0.337144), (58452,0.476549), (58453,0.353515), (58454,0.321990), (58455,0.225430), (58456,0.279370), (58457,0.227863), (58458,0.074172), (58459,0.511783), (58460,0.360878), (58461,0.258282), (58462,0.111561), (58463,0.375454), (58464,0.215257), (58465,0.183731), (58466,0.021675), (58467,0.572622), (58468,0.453771), (58469,0.413880), (58470,0.186802), (58471,0.557056), (58472,0.331838), (58473,0.169318), (58474,0.500562), (58475,0.360340), (58476,0.391982), (58477,0.252229), (58478,0.192826), (58479,0.049817), (58480,0.325790), (58481,0.200433), (58482,0.514482), (58483,0.355218), (58484,0.456534), (58485,0.298203), (58486,0.352136), (58487,0.228176), (58488,0.237989), (58489,0.055964), (58490,0.380239), (58491,0.239084), (58492,0.237752), (58493,0.068732), (58494,0.024658), (58495,-0.120668), (58496,0.026634), (58497,-0.129844), (58498,0.246453), (58499,0.064891), (58500,0.187108), (58501,0.030631), (58502,0.079924), (58503,-0.068657), (58504,0.058206), (58505,-0.080157), (58506,0.255734), (58507,0.110402), (58508,0.091875), (58509,-0.034872), (58510,-0.074300), (58511,-0.249819), (58512,0.029866), (58513,-0.123361), (58514,0.244576), (58515,0.090885), (58516,0.208919), (58517,0.039899), (58518,0.088266), (58519,-0.083540), (58520,0.244912), (58521,0.127451), (58522,0.100571), (58523,0.310576), (58524,0.309244), (58525,0.115604), (58526,0.082682), (58527,-0.109099), (58528,0.184055), (58529,-0.007262), (58530,-0.027179), (58531,0.171687), (58532,0.340817), (58533,0.190845), (58534,0.135162), (58535,0.094807), (58536,-0.146673), (58537,0.129293), (58538,0.370419), (58539,0.305913), (58540,0.173123), (58541,0.210338), (58542,0.008808), (58543,-0.051522), (58544,-0.180592), (58545,0.089332), (58546,0.322105), (58547,0.311944), (58548,0.133632), (58549,0.289292), (58550,0.226183), (58551,0.163993), (58552,-0.276751), (58553,0.018256), (58554,0.274248), (58555,0.154933), (58556,0.029576), (58557,0.026378), (58558,-0.089687), (58559,-0.140724), (58560,-0.328785), (58561,-0.000334), (58562,0.227793), (58563,0.157245), (58564,0.030028), (58565,0.156891), (58566,0.096104), (58567,0.022769), (58568,-0.175518), (58569,0.078157), (58570,0.311387), (58571,0.260350), (58572,0.121524), (58573,0.174067), (58574,-0.001452), (58575,-0.085006), (58576,-0.249843), (58577,0.025197), (58578,0.265859), (58579,0.188811), (58580,0.066704), (58581,0.175915), (58582,0.106300), (58583,0.091493), (58584,-0.057089), (58585,0.186360), (58586,0.084234), (58587,0.466104), (58588,0.295688), (58589,0.330586), (58590,0.110007), (58591,0.048288), (58592,-0.117019), (58593,0.164520), (58594,0.045206), (58595,0.349969), (58596,0.195352), (58597,0.353335), (58598,0.193602), (58599,0.249401), (58600,0.078985), (58601,0.324764), (58602,0.165963), (58603,0.531114), (58604,0.363484), (58605,0.373762), (58606,0.227966), (58607,0.147199), (58608,0.000477), (58609,0.285735), (58610,0.073053), (58611,0.444704), (58612,0.282653), (58613,0.414163), (58614,0.274404), (58615,0.298619), (58616,0.124027), (58617,0.429717), (58618,0.322938), (58619,0.642567), (58620,0.484699), (58621,0.434126), (58622,0.270679), (58623,0.170406), (58624,0.008356), (58625,0.306620), (58626,0.139923), (58627,0.449796), (58628,0.285422), (58629,0.460125), (58630,0.286929), (58631,0.314851), (58632,0.031568), (58633,0.307071), (58634,0.163599), (58635,0.485088), (58636,0.317928), (58637,0.319839), (58638,0.168934), (58639,0.089563), (58640,-0.056695), (58641,0.200229), (58642,0.049788), (58643,0.415865), (58644,0.200397), (58645,0.366276), (58646,0.193544), (58647,0.245160), (58648,0.206202), (58649,0.069229), (58650,0.050239), (58651,0.270470), (58652,0.276101), (58653,0.148884), (58654,0.101097), (58655,-0.087428), (58656,0.152772), (58657,0.015805), (58658,0.010748), (58659,0.252807), (58660,0.404291), (58661,0.265928), (58662,0.200489), (58663,0.122051), (58664,0.355281), (58665,0.235960), (58666,0.186783), (58667,0.418623), (58668,0.408925), (58669,0.198103), (58670,0.175863), (58671,-0.015918), (58672,0.277700), (58673,0.119362), (58674,0.083654), (58675,0.332682), (58676,0.492989), (58677,0.326292), (58678,0.255744), (58679,0.192634), (58680,0.354794), (58681,0.228047), (58682,0.175614), (58683,0.421392), (58684,0.447925), (58685,0.287264), (58686,0.194424), (58687,0.038873), (58688,0.330168), (58689,0.151856), (58690,0.143091), (58691,0.383291), (58692,0.498545), (58693,0.333238), (58694,0.299389), (58695,0.216298), (58696,0.398903), (58697,0.274009), (58698,0.196961), (58699,0.428338), (58700,0.450224), (58701,0.267272), (58702,0.233417), (58703,0.048142), (58704,0.340833), (58705,0.163917), (58706,0.074327), (58707,0.333105), (58708,0.522679), (58709,0.345763), (58710,0.308658), (58711,0.258547), (58712,0.334315), (58713,0.175984), (58714,0.123551), (58715,0.356318), (58716,0.372168), (58717,0.209190), (58718,0.117740), (58719,-0.031768), (58720,0.268813), (58721,0.092830), (58722,0.036214), (58723,0.292675), (58724,0.438580), (58725,0.292321), (58726,0.247790), (58727,0.163309), (58728,0.357523), (58729,0.162492), (58730,0.518814), (58731,0.374415), (58732,0.361468), (58733,0.215673), (58734,0.148374), (58735,-0.008104), (58736,0.266472), (58737,0.143902), (58738,0.455635), (58739,0.314949), (58740,0.430666), (58741,0.287658), (58742,0.292825), (58743,0.138671), (58744,0.185172), (58745,0.042169), (58746,0.380376), (58747,0.196955), (58748,0.187727), (58749,0.080948), (58750,0.004363), (58751,-0.166516), (58752,0.019802), (58753,-0.107409), (58754,0.236835), (58755,0.112874), (58756,0.220695), (58757,0.023342), (58758,0.082384), (58759,-0.070374), (58760,0.048130), (58761,-0.079550), (58762,0.308826), (58763,0.157458), (58764,0.142651), (58765,0.016361), (58766,-0.043499), (58767,-0.166533), (58768,0.084812), (58769,-0.059124), (58770,0.295809), (58771,0.138868), (58772,0.280126), (58773,0.110643), (58774,0.163656), (58775,0.001600), (58776,-0.025743), (58777,0.282270), (58778,0.124396), (58779,0.420337), (58780,0.271292), (58781,0.295971), (58782,0.193369), (58783,0.119107), (58784,-0.046193), (58785,0.232559), (58786,0.064936), (58787,0.450982), (58788,0.317266), (58789,0.449239), (58790,0.289975), (58791,0.336945), (58792,0.011390), (58793,0.267851), (58794,0.487612), (58795,0.408704), (58796,0.243867), (58797,0.239279), (58798,0.102313), (58799,0.035014), (58800,-0.139115), (58801,0.175868), (58802,0.410031), (58803,0.359927), (58804,0.184864), (58805,0.356323), (58806,0.235143), (58807,0.171100), (58808,-0.197185), (58809,0.083427), (58810,0.304585), (58811,0.263760), (58812,0.114716), (58813,0.142181), (58814,-0.036594), (58815,-0.090881), (58816,-0.276626), (58817,0.029534), (58818,0.259051), (58819,0.181076), (58820,0.037134), (58821,0.248073), (58822,0.136654), (58823,0.077721), (58824,-0.086659), (58825,0.168876), (58826,0.381204), (58827,0.345032), (58828,0.159288), (58829,0.193716), (58830,-0.009211), (58831,-0.049102), (58832,-0.221372), (58833,0.059704), (58834,0.324061), (58835,0.253976), (58836,0.110040), (58837,0.246659), (58838,0.204914), (58839,0.139475), (58840,-0.041154), (58841,0.238062), (58842,0.081585), (58843,0.419792), (58844,0.305587), (58845,0.308895), (58846,0.163563), (58847,0.101380), (58848,-0.065786), (58849,0.204144), (58850,0.028155), (58851,0.404452), (58852,0.197812), (58853,0.375307), (58854,0.195605), (58855,0.237466), (58856,0.064727), (58857,0.322114), (58858,0.192111), (58859,0.511276), (58860,0.361768), (58861,0.396660), (58862,0.266193), (58863,0.187285), (58864,0.040564), (58865,0.344400), (58866,0.153083), (58867,0.504302), (58868,0.343178), (58869,0.465858), (58870,0.358153), (58871,0.381436), (58872,0.240287), (58873,0.466554), (58874,0.322618), (58875,0.637138), (58876,0.457436), (58877,0.471426), (58878,0.360471), (58879,0.300604), (58880,0.076776), (58881,0.356456), (58882,0.186973), (58883,0.541905), (58884,0.368702), (58885,0.499748), (58886,0.330728), (58887,0.336823), (58888,0.024279), (58889,0.337865), (58890,0.217618), (58891,0.572550), (58892,0.377983), (58893,0.353890), (58894,0.217850), (58895,0.149625), (58896,0.007543), (58897,0.263077), (58898,0.088015), (58899,0.444343), (58900,0.292505), (58901,0.392894), (58902,0.274043), (58903,0.321477), (58904,0.391209), (58905,0.221726), (58906,0.159073), (58907,0.407168), (58908,0.398867), (58909,0.300917), (58910,0.281927), (58911,0.054380), (58912,0.354040), (58913,0.203599), (58914,0.134446), (58915,0.327270), (58916,0.488504), (58917,0.320880), (58918,0.318615), (58919,0.261999), (58920,0.390258), (58921,0.248646), (58922,0.165555), (58923,0.410401), (58924,0.428574), (58925,0.268847), (58926,0.194585), (58927,0.027888), (58928,0.322433), (58929,0.173851), (58930,0.106089), (58931,0.340715), (58932,0.505205), (58933,0.391927), (58934,0.336243), (58935,0.287993), (58936,0.432971), (58937,0.250482), (58938,0.221743), (58939,0.496313), (58940,0.494511), (58941,0.304590), (58942,0.276314), (58943,0.097538), (58944,0.392083), (58945,0.239325), (58946,0.172495), (58947,0.432670), (58948,0.528876), (58949,0.394690), (58950,0.340866), (58951,0.300048), (58952,0.455245), (58953,0.276476), (58954,0.226365), (58955,0.507441), (58956,0.546052), (58957,0.395611), (58958,0.368262), (58959,0.111453), (58960,0.404144), (58961,0.279714), (58962,0.242146), (58963,0.474919), (58964,0.580880), (58965,0.430902), (58966,0.408199), (58967,0.317682), (58968,0.490531), (58969,0.315006), (58970,0.303918), (58971,0.526466), (58972,0.552998), (58973,0.444359), (58974,0.368708), (58975,0.173214), (58976,0.509098), (58977,0.328469), (58978,0.309016), (58979,0.504626), (58980,0.635665), (58981,0.495913), (58982,0.430010), (58983,0.349243), (58984,0.406432), (58985,0.266679), (58986,0.623002), (58987,0.450269), (58988,0.472155), (58989,0.324970), (58990,0.189857), (58991,0.010618), (58992,0.280078), (58993,0.122674), (58994,0.441376), (58995,0.282576), (58996,0.446596), (58997,0.331927), (58998,0.417914), (58999,0.251218), (59000,0.237800), (59001,0.102694), (59002,0.426963), (59003,0.274205), (59004,0.329534), (59005,0.155405), (59006,0.043054), (59007,-0.132929), (59008,0.027841), (59009,-0.141179), (59010,0.245337), (59011,0.063312), (59012,0.234301), (59013,0.087116), (59014,0.136410), (59015,-0.020531), (59016,-0.193734), (59017,0.113816), (59018,0.386533), (59019,0.301588), (59020,0.141861), (59021,0.137736), (59022,-0.022461), (59023,-0.092076), (59024,-0.262486), (59025,0.018590), (59026,0.260179), (59027,0.189637), (59028,-0.001217), (59029,0.152590), (59030,0.121991), (59031,0.079776), (59032,-0.019107), (59033,0.240141), (59034,0.141728), (59035,0.452528), (59036,0.305806), (59037,0.309577), (59038,0.159136), (59039,0.080697), (59040,-0.070207), (59041,0.207149), (59042,0.069719), (59043,0.382842), (59044,0.237517), (59045,0.402470), (59046,0.291971), (59047,0.313394), (59048,-0.051641), (59049,0.213643), (59050,0.475677), (59051,0.443681), (59052,0.286277), (59053,0.251032), (59054,0.087585), (59055,-0.038699), (59056,-0.180311), (59057,0.130952), (59058,0.374871), (59059,0.348918), (59060,0.217518), (59061,0.367612), (59062,0.298454), (59063,0.207010), (59064,-0.264862), (59065,0.035725), (59066,0.281034), (59067,0.256008), (59068,0.124145), (59069,0.135819), (59070,-0.047603), (59071,-0.104213), (59072,-0.305280), (59073,-0.020491), (59074,0.222958), (59075,0.184926), (59076,0.045637), (59077,0.151599), (59078,0.096848), (59079,0.019330), (59080,-0.130178), (59081,0.133709), (59082,0.340465), (59083,0.303367), (59084,0.095794), (59085,0.152520), (59086,-0.002104), (59087,-0.077293), (59088,-0.207296), (59089,0.051488), (59090,0.312126), (59091,0.230431), (59092,0.082313), (59093,0.250053), (59094,0.177651), (59095,0.159587), (59096,-0.013146), (59097,0.234486), (59098,0.112843), (59099,0.484963), (59100,0.297365), (59101,0.316465), (59102,0.159524), (59103,0.102444), (59104,-0.058210), (59105,0.250736), (59106,0.074284), (59107,0.396699), (59108,0.256940), (59109,0.415394), (59110,0.222686), (59111,0.270583), (59112,0.117819), (59113,0.410973), (59114,0.231734), (59115,0.576447), (59116,0.411611), (59117,0.397730), (59118,0.248685), (59119,0.168381), (59120,0.058352), (59121,0.277657), (59122,0.152300), (59123,0.519304), (59124,0.411599), (59125,0.550077), (59126,0.361546), (59127,0.408517), (59128,0.193511), (59129,0.442540), (59130,0.346907), (59131,0.681401), (59132,0.521674), (59133,0.530091), (59134,0.368967), (59135,0.277054), (59136,0.041610), (59137,0.328265), (59138,0.176427), (59139,0.495593), (59140,0.384174), (59141,0.511501), (59142,0.343877), (59143,0.382489), (59144,0.100596), (59145,0.377952), (59146,0.236803), (59147,0.568511), (59148,0.443617), (59149,0.439962), (59150,0.250034), (59151,0.179956), (59152,0.055525), (59153,0.277146), (59154,0.162008), (59155,0.508581), (59156,0.384151), (59157,0.543994), (59158,0.391699), (59159,0.420091), (59160,0.400638), (59161,0.246020), (59162,0.205665), (59163,0.401739), (59164,0.412943), (59165,0.256928), (59166,0.186380), (59167,-0.001218), (59168,0.260816), (59169,0.142891), (59170,0.100213), (59171,0.345059), (59172,0.497470), (59173,0.324267), (59174,0.276016), (59175,0.209187), (59176,0.422449), (59177,0.284550), (59178,0.192636), (59179,0.464426), (59180,0.419888), (59181,0.278276), (59182,0.306668), (59183,0.108845), (59184,0.396890), (59185,0.250631), (59186,0.194948), (59187,0.436544), (59188,0.581985), (59189,0.418075), (59190,0.367038), (59191,0.301605), (59192,0.495355), (59193,0.341201), (59194,0.266933), (59195,0.538259), (59196,0.571761), (59197,0.375797), (59198,0.300145), (59199,0.149240), (59200,0.421950), (59201,0.237608), (59202,0.196784), (59203,0.438380), (59204,0.581968), (59205,0.443142), (59206,0.416719), (59207,0.355926), (59208,0.524129), (59209,0.314703), (59210,0.284104), (59211,0.504328), (59212,0.497417), (59213,0.339080), (59214,0.283403), (59215,0.135285), (59216,0.428902), (59217,0.271028), (59218,0.208382), (59219,0.447649), (59220,0.547574), (59221,0.379951), (59222,0.362820), (59223,0.302491), (59224,0.358284), (59225,0.178119), (59226,0.104790), (59227,0.351025), (59228,0.377558), (59229,0.245232), (59230,0.214169), (59231,0.002420), (59232,0.319262), (59233,0.174857), (59234,0.125679), (59235,0.357983), (59236,0.493205), (59237,0.350666), (59238,0.243888), (59239,0.238836), (59240,0.382418), (59241,0.241732), (59242,0.590165), (59243,0.443437), (59244,0.445818), (59245,0.262866), (59246,0.201146), (59247,0.044669), (59248,0.372194), (59249,0.193881), (59250,0.505614), (59251,0.348210), (59252,0.516876), (59253,0.341820), (59254,0.389717), (59255,0.235563), (59256,0.255126), (59257,0.085643), (59258,0.426179), (59259,0.269232), (59260,0.255358), (59261,0.123495), (59262,0.044587), (59263,-0.088666), (59264,0.237932), (59265,0.095857), (59266,0.011369), (59267,0.265971), (59268,0.429534), (59269,0.249831), (59270,0.166741), (59271,0.116167), (59272,0.003352), (59273,0.225436), (59274,0.070819), (59275,0.399740), (59276,0.288315), (59277,0.300445), (59278,0.129109), (59279,0.027440), (59280,-0.104887), (59281,0.196627), (59282,0.008102), (59283,0.336090), (59284,0.235354), (59285,0.372437), (59286,0.182515), (59287,0.248064), (59288,-0.051480), (59289,0.271868), (59290,0.152547), (59291,0.463353), (59292,0.333350), (59293,0.345017), (59294,0.185290), (59295,0.122637), (59296,-0.066814), (59297,0.208682), (59298,0.018761), (59299,0.356511), (59300,0.161944), (59301,0.369627), (59302,0.248452), (59303,0.261053), (59304,-0.201533), (59305,0.073506), (59306,0.275152), (59307,0.254309), (59308,0.123379), (59309,0.115072), (59310,-0.066484), (59311,-0.090120), (59312,-0.271682), (59313,0.045160), (59314,0.316023), (59315,0.274735), (59316,0.081564), (59317,0.220043), (59318,0.129056), (59319,0.097061), (59320,-0.058020), (59321,0.251853), (59322,0.022452), (59323,0.391779), (59324,0.220437), (59325,0.237213), (59326,0.095601), (59327,-0.020000), (59328,-0.108664), (59329,0.139901), (59330,-0.030978), (59331,0.304906), (59332,0.144252), (59333,0.281797), (59334,0.155977), (59335,0.156961), (59336,-0.057581), (59337,0.216532), (59338,0.091638), (59339,0.443321), (59340,0.285447), (59341,0.267853), (59342,0.135990), (59343,0.088672), (59344,-0.090566), (59345,0.197015), (59346,0.042391), (59347,0.377348), (59348,0.243169), (59349,0.395116), (59350,0.227950), (59351,0.250769), (59352,-0.062707), (59353,0.224405), (59354,0.096261), (59355,0.460485), (59356,0.315617), (59357,0.321248), (59358,0.171740), (59359,0.080290), (59360,-0.064572), (59361,0.177017), (59362,0.051197), (59363,0.351784), (59364,0.222244), (59365,0.365369), (59366,0.252084), (59367,0.253075), (59368,0.083122), (59369,0.348406), (59370,0.215616), (59371,0.595633), (59372,0.375054), (59373,0.410879), (59374,0.277156), (59375,0.223796), (59376,0.081257), (59377,0.316810), (59378,0.157546), (59379,0.533380), (59380,0.348105), (59381,0.502839), (59382,0.346361), (59383,0.379857), (59384,0.114689), (59385,0.379509), (59386,0.243470), (59387,0.571458), (59388,0.406621), (59389,0.429897), (59390,0.260884), (59391,0.170824), (59392,-0.194674), (59393,0.091974), (59394,-0.100270), (59395,0.278813), (59396,0.143243), (59397,0.287288), (59398,0.130348), (59399,0.158740), (59400,-0.211405), (59401,0.058055), (59402,-0.092380), (59403,0.269515), (59404,0.094923), (59405,0.139107), (59406,0.046267), (59407,-0.061439), (59408,-0.225349), (59409,0.033892), (59410,-0.093318), (59411,0.246279), (59412,0.100021), (59413,0.249181), (59414,0.115928), (59415,0.122956), (59416,0.295335), (59417,0.163478), (59418,0.039511), (59419,-0.079803), (59420,0.336437), (59421,0.210617), (59422,0.125672), (59423,-0.041951), (59424,0.188029), (59425,0.067319), (59426,-0.030637), (59427,-0.174573), (59428,0.396349), (59429,0.240335), (59430,0.179542), (59431,0.030961), (59432,0.272093), (59433,0.112829), (59434,0.074798), (59435,0.252756), (59436,0.225870), (59437,0.105622), (59438,0.023465), (59439,-0.147878), (59440,0.175933), (59441,0.053826), (59442,-0.003717), (59443,0.239275), (59444,0.374034), (59445,0.209198), (59446,0.155837), (59447,0.090398), (59448,0.136905), (59449,-0.004713), (59450,-0.056214), (59451,0.198387), (59452,0.195659), (59453,0.061943), (59454,0.037380), (59455,-0.172980), (59456,0.122492), (59457,-0.062320), (59458,-0.098955), (59459,0.144494), (59460,0.355432), (59461,0.190596), (59462,0.112151), (59463,0.037426), (59464,0.220030), (59465,0.033822), (59466,-0.040903), (59467,0.242496), (59468,0.246731), (59469,0.083753), (59470,0.022491), (59471,-0.121908), (59472,0.138730), (59473,-0.017285), (59474,-0.092010), (59475,0.157019), (59476,0.336367), (59477,0.154805), (59478,0.141395), (59479,0.054591), (59480,0.361214), (59481,0.209383), (59482,0.137907), (59483,-0.014857), (59484,0.405102), (59485,0.232370), (59486,0.122341), (59487,-0.001626), (59488,0.273877), (59489,0.127155), (59490,0.079368), (59491,-0.039484), (59492,0.474771), (59493,0.330829), (59494,0.230556), (59495,0.095913), (59496,0.137304), (59497,-0.003845), (59498,0.292560), (59499,0.197396), (59500,0.151932), (59501,-0.007332), (59502,-0.089953), (59503,-0.202768), (59504,0.075058), (59505,-0.081889), (59506,0.286512), (59507,0.161154), (59508,0.323321), (59509,0.166380), (59510,0.149250), (59511,-0.013727), (59512,0.221826), (59513,0.071385), (59514,0.021274), (59515,0.230359), (59516,0.254105), (59517,0.094372), (59518,0.044731), (59519,-0.088059), (59520,-0.018791), (59521,-0.144148), (59522,0.195919), (59523,0.005528), (59524,0.175591), (59525,0.038161), (59526,0.071657), (59527,-0.069956), (59528,-0.259413), (59529,0.009590), (59530,0.237247), (59531,0.184350), (59532,0.005111), (59533,0.040473), (59534,-0.164777), (59535,-0.208382), (59536,-0.357433), (59537,-0.094936), (59538,0.158739), (59539,0.154151), (59540,-0.038557), (59541,0.114781), (59542,0.044232), (59543,-0.013768), (59544,-0.376950), (59545,-0.091691), (59546,0.139216), (59547,0.074710), (59548,-0.088274), (59549,-0.009713), (59550,-0.228901), (59551,-0.290621), (59552,-0.463817), (59553,-0.183675), (59554,0.076500), (59555,0.031505), (59556,-0.155166), (59557,0.031615), (59558,-0.075627), (59559,-0.102507), (59560,-0.289642), (59561,0.034627), (59562,0.260894), (59563,0.208467), (59564,0.028295), (59565,0.032073), (59566,-0.151812), (59567,-0.224684), (59568,-0.343072), (59569,-0.081971), (59570,0.175417), (59571,0.102551), (59572,-0.054396), (59573,0.119386), (59574,0.058593), (59575,-0.024028), (59576,-0.374667), (59577,-0.126109), (59578,0.141961), (59579,0.062590), (59580,-0.112929), (59581,-0.084074), (59582,-0.211754), (59583,-0.195441), (59584,-0.361204), (59585,-0.134010), (59586,0.149852), (59587,0.127149), (59588,-0.059986), (59589,0.101711), (59590,0.049284), (59591,-0.037520), (59592,-0.231161), (59593,0.044805), (59594,0.350502), (59595,0.268807), (59596,0.116513), (59597,0.158837), (59598,-0.063138), (59599,-0.156905), (59600,-0.291091), (59601,-0.063427), (59602,0.179559), (59603,0.114120), (59604,-0.006591), (59605,0.141173), (59606,0.071095), (59607,0.006119), (59608,-0.391897), (59609,-0.047647), (59610,0.172114), (59611,0.127583), (59612,-0.087422), (59613,-0.007472), (59614,-0.187174), (59615,-0.250753), (59616,-0.406767), (59617,-0.132198), (59618,0.107539), (59619,0.078336), (59620,-0.140852), (59621,0.055221), (59622,-0.029723), (59623,-0.105845), (59624,-0.249317), (59625,0.013644), (59626,0.234802), (59627,0.161467), (59628,0.050975), (59629,0.056142), (59630,-0.159326), (59631,-0.161592), (59632,-0.306923), (59633,-0.059755), (59634,0.187414), (59635,0.153095), (59636,0.011946), (59637,0.158321), (59638,0.076163), (59639,-0.010177), (59640,-0.105341), (59641,0.191064), (59642,0.031336), (59643,0.354678), (59644,0.218639), (59645,0.201045), (59646,0.062219), (59647,0.022328), (59648,-0.136473), (59649,0.153432), (59650,0.002991), (59651,0.332838), (59652,0.205158), (59653,0.345490), (59654,0.160215), (59655,0.128220), (59656,-0.154136), (59657,0.135768), (59658,0.035959), (59659,0.373239), (59660,0.193074), (59661,0.213100), (59662,0.061732), (59663,-0.007420), (59664,-0.153215), (59665,0.090234), (59666,-0.035586), (59667,0.308200), (59668,0.200025), (59669,0.305523), (59670,0.134650), (59671,0.170469), (59672,0.231378), (59673,0.073967), (59674,-0.004008), (59675,0.253843), (59676,0.231604), (59677,0.087668), (59678,0.048703), (59679,-0.106378), (59680,0.168198), (59681,0.041908), (59682,-0.065334), (59683,0.171616), (59684,0.343538), (59685,0.176841), (59686,0.119762), (59687,0.058505), (59688,0.089221), (59689,-0.038460), (59690,0.296034), (59691,0.094034), (59692,0.119640), (59693,-0.021509), (59694,-0.125501), (59695,-0.232743), (59696,0.031151), (59697,-0.143912), (59698,0.216593), (59699,0.038751), (59700,0.157718), (59701,0.018892), (59702,0.061217), (59703,-0.093865), (59704,0.182101), (59705,0.060921), (59706,0.001061), (59707,0.212926), (59708,0.221807), (59709,0.071835), (59710,0.017542), (59711,-0.168196), (59712,0.131458), (59713,0.007034), (59714,-0.064442), (59715,0.192946), (59716,0.357429), (59717,0.160076), (59718,0.144342), (59719,0.082159), (59720,0.258721), (59721,0.115712), (59722,0.067461), (59723,0.275614), (59724,0.318871), (59725,0.139632), (59726,0.096021), (59727,-0.061383), (59728,0.199254), (59729,0.062752), (59730,0.021470), (59731,0.251914), (59732,0.372277), (59733,0.262712), (59734,0.187054), (59735,0.127194), (59736,0.289354), (59737,0.181649), (59738,0.117143), (59739,0.351770), (59740,0.336962), (59741,0.191631), (59742,0.149886), (59743,-0.097167), (59744,0.208060), (59745,0.033931), (59746,-0.003638), (59747,0.231922), (59748,0.406624), (59749,0.242251), (59750,0.248815), (59751,0.163864), (59752,-0.085048), (59753,0.188131), (59754,0.437623), (59755,0.392159), (59756,0.251473), (59757,0.233416), (59758,0.063470), (59759,-0.016365), (59760,-0.148691), (59761,0.126348), (59762,0.302910), (59763,0.282067), (59764,0.128376), (59765,0.314230), (59766,0.176794), (59767,0.173603), (59768,0.226146), (59769,0.049230), (59770,0.398120), (59771,0.227710), (59772,0.227768), (59773,0.082900), (59774,-0.008081), (59775,-0.107427), (59776,0.008754), (59777,-0.173735), (59778,0.188160), (59779,0.059090), (59780,0.202672), (59781,0.062450), (59782,0.046716), (59783,-0.113011), (59784,0.070983), (59785,-0.093390), (59786,0.209520), (59787,0.059078), (59788,0.078642), (59789,-0.029990), (59790,-0.134446), (59791,-0.264449), (59792,0.036138), (59793,-0.117090), (59794,0.189997), (59795,0.057677), (59796,0.165028), (59797,0.059183), (59798,0.045766), (59799,-0.073085), (59800,-0.399567), (59801,-0.125461), (59802,0.135176), (59803,0.047909), (59804,-0.118324), (59805,-0.074603), (59806,-0.244550), (59807,-0.287691), (59808,-0.438132), (59809,-0.142655), (59810,0.093825), (59811,0.027459), (59812,-0.159675), (59813,-0.017947), (59814,-0.073630), (59815,-0.112589), (59816,-0.325735), (59817,-0.056738), (59818,0.229917), (59819,0.178874), (59820,-0.001292), (59821,-0.004020), (59822,-0.169790), (59823,-0.205962), (59824,-0.345721), (59825,-0.066035), (59826,0.227119), (59827,0.155180), (59828,-0.018949), (59829,0.107914), (59830,0.063840), (59831,0.006766), (59832,-0.367561), (59833,-0.041890), (59834,0.223857), (59835,0.180716), (59836,0.020519), (59837,-0.007294), (59838,-0.142870), (59839,-0.191120), (59840,-0.381505), (59841,-0.082778), (59842,0.153709), (59843,0.078514), (59844,-0.106298), (59845,0.041003), (59846,-0.029539), (59847,-0.040170), (59848,-0.221731), (59849,0.088148), (59850,0.301403), (59851,0.269878), (59852,0.127332), (59853,0.119031), (59854,-0.078323), (59855,-0.167450), (59856,-0.290484), (59857,0.004524), (59858,0.235901), (59859,0.189046), (59860,0.020953), (59861,0.154322), (59862,0.074018), (59863,0.007189), (59864,-0.383394), (59865,-0.126469), (59866,0.130449), (59867,0.107282), (59868,-0.038050), (59869,-0.063539), (59870,-0.222803), (59871,-0.279877), (59872,-0.463298), (59873,-0.170607), (59874,0.097463), (59875,0.047353), (59876,-0.091473), (59877,0.042359), (59878,-0.051414), (59879,-0.053679), (59880,-0.233845), (59881,0.004958), (59882,0.270242), (59883,0.213632), (59884,0.007919), (59885,0.001471), (59886,-0.119703), (59887,-0.170277), (59888,-0.314212), (59889,-0.032210), (59890,0.213569), (59891,0.166708), (59892,-0.005562), (59893,0.153818), (59894,0.043320), (59895,-0.023972), (59896,-0.090801), (59897,0.208853), (59898,0.083959), (59899,0.406844), (59900,0.267085), (59901,0.286654), (59902,0.152005), (59903,0.048946), (59904,-0.114038), (59905,0.168898), (59906,0.031925), (59907,0.355737), (59908,0.209478), (59909,0.374431), (59910,0.234672), (59911,0.257491), (59912,-0.079673), (59913,0.191647), (59914,0.037493), (59915,0.394748), (59916,0.264281), (59917,0.222993), (59918,0.063266), (59919,0.009906), (59920,-0.114988), (59921,0.134504), (59922,-0.068423), (59923,0.318556), (59924,0.182517), (59925,0.313563), (59926,0.177060), (59927,0.228207), (59928,0.261709), (59929,0.072714), (59930,0.043975), (59931,0.291144), (59932,0.274477), (59933,0.138901), (59934,0.074858), (59935,-0.090912), (59936,0.159513), (59937,-0.016013), (59938,-0.065190), (59939,0.176399), (59940,0.367363), (59941,0.207172), (59942,0.168677), (59943,0.106488), (59944,0.128381), (59945,-0.056431), (59946,0.266911), (59947,0.132731), (59948,0.137429), (59949,0.000463), (59950,-0.075659), (59951,-0.233063), (59952,0.048476), (59953,-0.099642), (59954,0.202335), (59955,0.016597), (59956,0.173184), (59957,0.038077), (59958,0.068323), (59959,-0.055638), (59960,0.244480), (59961,0.096831), (59962,0.038825), (59963,0.272055), (59964,0.291624), (59965,0.085911), (59966,0.042770), (59967,-0.155517), (59968,0.139497), (59969,-0.016054), (59970,-0.062445), (59971,0.181468), (59972,0.380797), (59973,0.230820), (59974,0.188611), (59975,0.079510), (59976,0.277906), (59977,0.110276), (59978,0.077824), (59979,0.323596), (59980,0.329690), (59981,0.179719), (59982,0.088269), (59983,-0.091433), (59984,0.196612), (59985,-0.005388), (59986,0.006742), (59987,0.283178), (59988,0.393779), (59989,0.277251), (59990,0.216922), (59991,0.128728), (59992,0.290888), (59993,0.153458), (59994,0.086629), (59995,0.321719), (59996,0.344532), (59997,0.221498), (59998,0.132371), (59999,-0.036179), (60000,0.253719), (60001,0.058689), (60002,0.006262), (60003,0.235309), (60004,0.416987), (60005,0.237748), (60006,0.211795), (60007,0.168654), (60008,0.193790), (60009,0.074006), (60010,0.384812), (60011,0.202323), (60012,0.243257), (60013,0.087707), (60014,0.039456), (60015,-0.123064), (60016,0.160334), (60017,-0.016581), (60018,0.314663), (60019,0.156326), (60020,0.321742), (60021,0.165264), (60022,0.157426), (60023,0.033466), (60024,0.122239), (60025,-0.039348), (60026,0.259379), (60027,0.105225), (60028,0.100637), (60029,-0.069316), (60030,-0.111524), (60031,-0.272184), (60032,-0.438418), (60033,-0.181493), (60034,0.089363), (60035,0.082915), (60036,-0.081458), (60037,0.113689), (60038,0.013879), (60039,-0.044591), (60040,-0.336239), (60041,-0.018933), (60042,0.217553), (60043,0.186027), (60044,0.024903), (60045,0.009633), (60046,-0.166819), (60047,-0.185809), (60048,-0.365048), (60049,-0.071430), (60050,0.150654), (60051,0.120518), (60052,-0.072653), (60053,0.073722), (60054,-0.029807), (60055,-0.051114), (60056,-0.194586), (60057,-0.319480), (60058,0.334585), (60059,0.201795), (60060,0.137289), (60061,-0.018725), (60062,0.005021), (60063,-0.140311), (60064,-0.195061), (60065,-0.359434), (60066,0.318781), (60067,0.147908), (60068,0.114053), (60069,-0.072149), (60070,0.133674), (60071,0.032475), (60072,-0.308872), (60073,-0.090038), (60074,0.198934), (60075,0.046633), (60076,0.009534), (60077,-0.167382), (60078,-0.182652), (60079,-0.333557), (60080,-0.369735), (60081,-0.103982), (60082,0.160369), (60083,0.016434), (60084,-0.055042), (60085,-0.146029), (60086,0.036576), (60087,-0.134303), (60088,-0.250831), (60089,-0.367829), (60090,0.294132), (60091,0.165988), (60092,0.122383), (60093,-0.074037), (60094,-0.080949), (60095,-0.236499), (60096,-0.304262), (60097,-0.437515), (60098,0.221660), (60099,0.058219), (60100,0.000213), (60101,-0.159984), (60102,0.080685), (60103,-0.090195), (60104,-0.217411), (60105,-0.321397), (60106,0.368897), (60107,0.208700), (60108,0.163242), (60109,0.001655), (60110,0.013786), (60111,-0.157557), (60112,-0.170504), (60113,-0.378541), (60114,0.315467), (60115,0.185007), (60116,0.126537), (60117,-0.030410), (60118,0.159627), (60119,0.034734), (60120,-0.152401), (60121,-0.283794), (60122,0.405110), (60123,0.276497), (60124,0.192480), (60125,-0.002081), (60126,0.004476), (60127,-0.159897), (60128,-0.207685), (60129,-0.365089), (60130,0.323809), (60131,0.160832), (60132,0.117221), (60133,-0.038323), (60134,0.203736), (60135,0.027284), (60136,-0.057197), (60137,-0.176981), (60138,0.501235), (60139,0.332685), (60140,0.298366), (60141,0.127023), (60142,0.130331), (60143,-0.021964), (60144,-0.060922), (60145,-0.229015), (60146,0.467322), (60147,0.316418), (60148,0.217535), (60149,0.039693), (60150,0.295221), (60151,0.129914), (60152,-0.087878), (60153,-0.249465), (60154,0.461268), (60155,0.308510), (60156,0.246321), (60157,0.059656), (60158,0.035556), (60159,-0.093051), (60160,-0.099035), (60161,-0.339582), (60162,0.359999), (60163,0.201198), (60164,0.154807), (60165,-0.010493), (60166,0.213914), (60167,0.089021), (60168,-0.160818), (60169,-0.280603), (60170,0.346518), (60171,0.246245), (60172,0.154795), (60173,-0.004932), (60174,0.003022), (60175,-0.168321), (60176,-0.224004), (60177,-0.349825), (60178,0.331184), (60179,0.183993), (60180,0.074897), (60181,-0.048607), (60182,0.210178), (60183,0.097363), (60184,-0.190103), (60185,0.063102), (60186,0.314447), (60187,0.274099), (60188,0.093927), (60189,0.091199), (60190,-0.105228), (60191,-0.164162), (60192,-0.304378), (60193,0.000849), (60194,0.239659), (60195,0.210913), (60196,0.028888), (60197,0.170153), (60198,0.120042), (60199,0.047640), (60200,-0.152037), (60201,0.129502), (60202,0.383177), (60203,0.360004), (60204,0.205386), (60205,0.170604), (60206,-0.014671), (60207,-0.074530), (60208,-0.192455), (60209,0.079328), (60210,0.307919), (60211,0.252235), (60212,0.094361), (60213,0.224944), (60214,0.167864), (60215,0.136802), (60216,-0.185497), (60217,0.100218), (60218,0.351570), (60219,0.274985), (60220,0.107361), (60221,0.127851), (60222,-0.034663), (60223,-0.101492), (60224,-0.239391), (60225,0.022643), (60226,0.258196), (60227,0.206226), (60228,0.082265), (60229,0.263474), (60230,0.154842), (60231,0.092189), (60232,-0.194344), (60233,0.089982), (60234,0.304634), (60235,0.277754), (60236,0.113844), (60237,0.133407), (60238,-0.012388), (60239,-0.076431), (60240,-0.225939), (60241,0.024943), (60242,0.286977), (60243,0.239652), (60244,0.046012), (60245,0.243482), (60246,0.140422), (60247,0.128402), (60248,-0.129803), (60249,0.130371), (60250,0.332950), (60251,0.326503), (60252,0.161202), (60253,0.181229), (60254,-0.038886), (60255,-0.082954), (60256,-0.206451), (60257,0.080660), (60258,0.366846), (60259,0.279578), (60260,0.137033), (60261,0.244391), (60262,0.193817), (60263,0.166931), (60264,-0.229688), (60265,0.457821), (60266,0.302739), (60267,0.242873), (60268,0.099401), (60269,0.093417), (60270,-0.057482), (60271,-0.107129), (60272,-0.297977), (60273,0.353765), (60274,0.194501), (60275,0.131848), (60276,-0.038561), (60277,0.209534), (60278,0.063739), (60279,0.002946), (60280,-0.174433), (60281,0.135440), (60282,0.401650), (60283,0.319493), (60284,0.174630), (60285,0.211382), (60286,0.033533), (60287,-0.037942), (60288,-0.326798), (60289,-0.470270), (60290,0.218165), (60291,0.036610), (60292,-0.054840), (60293,-0.240585), (60294,-0.005958), (60295,-0.130846), (60296,-0.269678), (60297,-0.434515), (60298,0.271108), (60299,0.104875), (60300,0.045479), (60301,-0.131437), (60302,-0.126733), (60303,-0.278101), (60304,-0.299414), (60305,-0.447062), (60306,0.174949), (60307,0.018471), (60308,-0.006092), (60309,-0.176965), (60310,0.051156), (60311,-0.098352), (60312,-0.115019), (60313,-0.297045), (60314,-0.047553), (60315,0.249315), (60316,0.176913), (60317,0.016252), (60318,0.028389), (60319,-0.142954), (60320,-0.193064), (60321,-0.348152), (60322,-0.094477), (60323,0.121571), (60324,0.083539), (60325,-0.086413), (60326,0.052992), (60327,-0.050067), (60328,-0.222800), (60329,-0.356986), (60330,0.318913), (60331,0.152217), (60332,0.069596), (60333,-0.071090), (60334,-0.101226), (60335,-0.243771), (60336,-0.276230), (60337,-0.438744), (60338,0.304036), (60339,0.158711), (60340,0.053322), (60341,-0.092936), (60342,0.114289), (60343,0.025162), (60344,-0.330587), (60345,-0.481955), (60346,0.200914), (60347,0.013309), (60348,-0.032619), (60349,-0.157043), (60350,-0.183465), (60351,-0.335297), (60352,-0.407235), (60353,-0.557677), (60354,0.098248), (60355,-0.026646), (60356,-0.106480), (60357,-0.227655), (60358,-0.006967), (60359,-0.177376), (60360,-0.203336), (60361,-0.380251), (60362,0.251985), (60363,0.124768), (60364,0.095566), (60365,-0.071131), (60366,-0.053428), (60367,-0.242885), (60368,-0.270698), (60369,-0.453186), (60370,0.210171), (60371,0.115934), (60372,0.032850), (60373,-0.100403), (60374,0.148619), (60375,-0.019005), (60376,-0.122997), (60377,-0.329637), (60378,0.005321), (60379,0.196285), (60380,0.169399), (60381,0.024530), (60382,0.050136), (60383,-0.115164), (60384,-0.207078), (60385,-0.405828), (60386,-0.105704), (60387,0.157256), (60388,0.089958), (60389,-0.088812), (60390,0.074282), (60391,0.039963), (60392,-0.006428), (60393,-0.085799), (60394,-0.217662), (60395,0.467993), (60396,0.317551), (60397,0.270227), (60398,0.094245), (60399,0.046457), (60400,-0.102124), (60401,-0.119718), (60402,-0.283165), (60403,0.410386), (60404,0.278986), (60405,0.205188), (60406,-0.031182), (60407,0.233175), (60408,0.040004), (60409,-0.124376), (60410,0.165065), (60411,0.398295), (60412,0.369556), (60413,0.195890), (60414,0.239148), (60415,0.039471), (60416,0.018621), (60417,-0.109523), (60418,0.160871), (60419,0.357414), (60420,0.253422), (60421,0.124345), (60422,0.265147), (60423,0.221079), (60424,-0.005072), (60425,-0.050073), (60426,-0.202838), (60427,0.487927), (60428,0.327730), (60429,0.278089), (60430,0.132294), (60431,0.124919), (60432,-0.017626), (60433,-0.035220), (60434,-0.187521), (60435,0.470727), (60436,0.306816), (60437,0.203294), (60438,0.073754), (60439,0.320459), (60440,-0.059441), (60441,0.235103), (60442,0.093028), (60443,0.449813), (60444,0.261289), (60445,0.296644), (60446,0.127161), (60447,0.047789), (60448,-0.089647), (60449,0.171461), (60450,0.027056), (60451,0.371305), (60452,0.206932), (60453,0.358416), (60454,0.193573), (60455,0.253549), (60456,0.068737), (60457,-0.116075), (60458,0.183579), (60459,0.427035), (60460,0.344877), (60461,0.187936), (60462,0.215395), (60463,0.064491), (60464,0.028319), (60465,-0.129555), (60466,0.144557), (60467,0.376391), (60468,0.352761), (60469,0.196747), (60470,0.325470), (60471,0.254458), (60472,-0.024648), (60473,0.259684), (60474,0.124108), (60475,0.485076), (60476,0.316056), (60477,0.359777), (60478,0.202366), (60479,0.083979), (60480,-0.077145), (60481,0.154232), (60482,0.027948), (60483,0.354539), (60484,0.214787), (60485,0.339790), (60486,0.198178), (60487,0.194053), (60488,0.028753), (60489,-0.087318), (60490,0.164497), (60491,0.436750), (60492,0.431229), (60493,0.237594), (60494,0.235329), (60495,0.085815), (60496,-0.006562), (60497,-0.148174), (60498,0.156126), (60499,0.368924), (60500,0.325783), (60501,0.168372), (60502,0.293382), (60503,0.287398), (60504,-0.000995), (60505,0.268002), (60506,0.118494), (60507,0.423721), (60508,0.289078), (60509,0.301672), (60510,0.174924), (60511,0.086724), (60512,-0.060461), (60513,0.180665), (60514,0.018615), (60515,0.371687), (60516,0.219392), (60517,0.342073), (60518,0.213466), (60519,0.261833), (60520,-0.012164), (60521,-0.154246), (60522,0.465448), (60523,0.349847), (60524,0.350832), (60525,0.210610), (60526,0.202772), (60527,0.011460), (60528,-0.060015), (60529,-0.198847), (60530,0.480765), (60531,0.306636), (60532,0.267214), (60533,0.088902), (60534,0.317029), (60535,0.121065), (60536,-0.217959), (60537,-0.348425), (60538,0.336766), (60539,0.193294), (60540,0.110204), (60541,0.004358), (60542,-0.014169), (60543,-0.147885), (60544,-0.384719), (60545,-0.531440), (60546,0.151422), (60547,0.032101), (60548,-0.006858), (60549,-0.148940), (60550,0.099625), (60551,-0.062895), (60552,-0.265821), (60553,-0.396751), (60554,0.225266), (60555,0.057637), (60556,0.022398), (60557,-0.147555), (60558,-0.162826), (60559,-0.310011), (60560,-0.349439), (60561,-0.521708), (60562,0.133283), (60563,-0.026908), (60564,-0.080268), (60565,-0.204235), (60566,-0.021167), (60567,-0.149310), (60568,-0.192452), (60569,-0.325705), (60570,-0.035337), (60571,0.130079), (60572,0.112949), (60573,-0.049565), (60574,-0.026752), (60575,-0.218063), (60576,-0.255631), (60577,-0.439046), (60578,-0.129173), (60579,0.110099), (60580,0.096682), (60581,-0.085343), (60582,0.055922), (60583,-0.029955), (60584,-0.248210), (60585,-0.420943), (60586,0.253560), (60587,0.124020), (60588,0.047435), (60589,-0.093714), (60590,-0.147538), (60591,-0.271968), (60592,-0.301171), (60593,-0.476227), (60594,0.173192), (60595,0.038079), (60596,-0.015745), (60597,-0.215421), (60598,0.043363), (60599,-0.034619), (60600,-0.340199), (60601,-0.535230), (60602,0.165284), (60603,-0.024637), (60604,-0.094716), (60605,-0.246090), (60606,-0.243246), (60607,-0.366280), (60608,-0.423817), (60609,-0.584940), (60610,0.092349), (60611,-0.124047), (60612,-0.130031), (60613,-0.282796), (60614,-0.083003), (60615,-0.249236), (60616,-0.322101), (60617,-0.504126), (60618,0.192204), (60619,0.053379), (60620,0.006988), (60621,-0.173184), (60622,-0.157334), (60623,-0.322171), (60624,-0.380178), (60625,-0.511571), (60626,0.162469), (60627,0.035252), (60628,-0.025541), (60629,-0.205243), (60630,0.043322), (60631,-0.088541), (60632,-0.182778), (60633,-0.336469), (60634,-0.039601), (60635,0.227079), (60636,0.139812), (60637,-0.008307), (60638,-0.010572), (60639,-0.179128), (60640,-0.219946), (60641,-0.385246), (60642,-0.111140), (60643,0.141602), (60644,0.089168), (60645,-0.069163), (60646,0.053517), (60647,0.007590), (60648,-0.032765), (60649,-0.128861), (60650,-0.289515), (60651,0.399383), (60652,0.251734), (60653,0.170967), (60654,0.031214), (60655,0.050314), (60656,-0.132175), (60657,-0.173926), (60658,-0.298820), (60659,0.352928), (60660,0.186232), (60661,0.133335), (60662,-0.009674), (60663,0.202655), (60664,-0.012814), (60665,-0.132592), (60666,0.132686), (60667,0.404475), (60668,0.327427), (60669,0.156548), (60670,0.205841), (60671,-0.022633), (60672,-0.025362), (60673,-0.189272), (60674,0.104346), (60675,0.368233), (60676,0.300008), (60677,0.123562), (60678,0.318702), (60679,0.253733), (60680,0.063342), (60681,-0.026712), (60682,-0.159032), (60683,0.467626), (60684,0.367816), (60685,0.296804), (60686,0.161692), (60687,0.150141), (60688,-0.031885), (60689,-0.071776), (60690,-0.228254), (60691,0.416519), (60692,0.240536), (60693,0.205754), (60694,0.068318), (60695,0.301555), (60696,-0.198188), (60697,0.106582), (60698,-0.056401), (60699,0.302244), (60700,0.117896), (60701,0.145361), (60702,-0.019482), (60703,-0.126718), (60704,-0.245112), (60705,0.006703), (60706,-0.161853), (60707,0.205621), (60708,0.058429), (60709,0.218273), (60710,0.068764), (60711,0.087864), (60712,-0.020768), (60713,-0.195824), (60714,0.082465), (60715,0.369577), (60716,0.342228), (60717,0.139765), (60718,0.147719), (60719,-0.032910), (60720,-0.077448), (60721,-0.233925), (60722,0.066662), (60723,0.315684), (60724,0.292517), (60725,0.129070), (60726,0.258720), (60727,0.169599), (60728,-0.081636), (60729,0.200366), (60730,0.004872), (60731,0.360731), (60732,0.200540), (60733,0.218244), (60734,0.035755), (60735,-0.068237), (60736,-0.225178), (60737,0.056831), (60738,-0.019291), (60739,0.310094), (60740,0.174518), (60741,0.282802), (60742,0.099844), (60743,0.128236), (60744,-0.044497), (60745,-0.182396), (60746,0.117722), (60747,0.445246), (60748,0.385850), (60749,0.247487), (60750,0.209456), (60751,0.058551), (60752,0.007977), (60753,-0.171725), (60754,0.119570), (60755,0.330045), (60756,0.287830), (60757,0.114171), (60758,0.264722), (60759,0.200216), (60760,-0.149960), (60761,0.106031), (60762,-0.032795), (60763,0.354191), (60764,0.197707), (60765,0.190802), (60766,0.045933), (60767,-0.018109), (60768,-0.138820), (60769,0.099983), (60770,-0.077859), (60771,0.233410), (60772,0.119662), (60773,0.292048), (60774,0.096554), (60775,0.103575), (60776,-0.058013), (60777,-0.181046), (60778,0.479987), (60779,0.357880), (60780,0.303593), (60781,0.135507), (60782,0.133705), (60783,-0.019060), (60784,-0.092858), (60785,-0.218678), (60786,0.429813), (60787,0.254758), (60788,0.176313), (60789,0.041200), (60790,0.251212), (60791,0.121209), (60792,-0.164397), (60793,-0.346422), (60794,0.324825), (60795,0.192041), (60796,0.159583), (60797,0.035152), (60798,-0.004270), (60799,-0.146815), (60800,-0.199712), (60801,-0.399389), (60802,-0.167085), (60803,0.131179), (60804,0.123804), (60805,-0.023851), (60806,0.115555), (60807,0.035720), (60808,-0.131440), (60809,-0.314392), (60810,-0.035176), (60811,0.215706), (60812,0.173961), (60813,-0.002955), (60814,0.023114), (60815,-0.160771), (60816,-0.193229), (60817,-0.326019), (60818,-0.051906), (60819,0.193403), (60820,0.119141), (60821,-0.036873), (60822,0.102995), (60823,-0.008423), (60824,-0.226685), (60825,-0.378053), (60826,-0.096508), (60827,0.125577), (60828,0.075466), (60829,-0.076365), (60830,-0.058192), (60831,-0.243004), (60832,-0.258744), (60833,-0.384564), (60834,-0.163407), (60835,0.092585), (60836,0.051767), (60837,-0.091705), (60838,0.056992), (60839,0.004559), (60840,-0.101287), (60841,-0.287495), (60842,-0.000846), (60843,0.243536), (60844,0.160915), (60845,0.002577), (60846,0.030506), (60847,-0.145483), (60848,-0.190020), (60849,-0.325127), (60850,-0.026400), (60851,0.170601), (60852,0.110741), (60853,-0.063858), (60854,0.090412), (60855,0.034729), (60856,-0.158442), (60857,-0.316779), (60858,-0.079830), (60859,0.186381), (60860,0.106546), (60861,-0.027170), (60862,-0.041977), (60863,-0.229112), (60864,-0.245779), (60865,-0.419908), (60866,-0.181562), (60867,0.069783), (60868,0.061482), (60869,-0.107538), (60870,0.021648), (60871,-0.020097), (60872,-0.079036), (60873,-0.211820), (60874,0.090158), (60875,0.311315), (60876,0.257485), (60877,0.096831), (60878,0.115004), (60879,-0.039620), (60880,-0.111095), (60881,-0.314485), (60882,-0.028300), (60883,0.189138), (60884,0.189196), (60885,0.026219), (60886,0.174447), (60887,0.103435), (60888,-0.216547), (60889,-0.341435), (60890,-0.047354), (60891,0.196096), (60892,0.112548), (60893,-0.050436), (60894,-0.036445), (60895,-0.175735), (60896,-0.259752), (60897,-0.405547), (60898,-0.094278), (60899,0.094826), (60900,0.009419), (60901,-0.111292), (60902,0.058764), (60903,0.001227), (60904,-0.063748), (60905,-0.122682), (60906,-0.333504), (60907,0.360047), (60908,0.224001), (60909,0.167391), (60910,0.001157), (60911,0.024903), (60912,-0.155262), (60913,-0.195617), (60914,-0.372532), (60915,0.296861), (60916,0.161285), (60917,0.113967), (60918,-0.019756), (60919,0.212554), (60920,0.018450), (60921,-0.140351), (60922,0.105885), (60923,0.382321), (60924,0.338247), (60925,0.161801), (60926,0.145134), (60927,-0.054543), (60928,-0.124622), (60929,-0.282496), (60930,0.016231), (60931,0.263400), (60932,0.203997), (60933,0.064245), (60934,0.194357), (60935,0.110810), (60936,-0.082831), (60937,-0.119936), (60938,-0.297778), (60939,0.388340), (60940,0.256940), (60941,0.200794), (60942,0.042926), (60943,0.003498), (60944,-0.102811), (60945,-0.177543), (60946,-0.342379), (60947,0.358134), (60948,0.166817), (60949,0.165021), (60950,0.031768), (60951,0.218086), (60952,-0.039655), (60953,0.242817), (60954,0.123496), (60955,0.036692), (60956,0.272715), (60957,0.263944), (60958,0.114899), (60959,0.042034), (60960,-0.097725), (60961,0.200539), (60962,0.004575), (60963,-0.072010), (60964,0.160763), (60965,0.321533), (60966,0.167842), (60967,0.102403), (60968,-0.150222), (60969,-0.325278), (60970,-0.033983), (60971,0.223398), (60972,0.206274), (60973,-0.005945), (60974,-0.004960), (60975,-0.198131), (60976,-0.207366), (60977,-0.397287), (60978,-0.097169), (60979,0.202491), (60980,0.110578), (60981,-0.047296), (60982,0.108834), (60983,0.083808), (60984,-0.211554), (60985,0.104819), (60986,-0.061878), (60987,0.258684), (60988,0.116139), (60989,0.121770), (60990,-0.064902), (60991,-0.155882), (60992,-0.293318), (60993,0.000300), (60994,-0.165933), (60995,0.192712), (60996,0.055282), (60997,0.164957), (60998,0.056788), (60999,0.035945), (61000,-0.098241), (61001,-0.306741), (61002,-0.040994), (61003,0.184341), (61004,0.168143), (61005,0.007483), (61006,0.026119), (61007,-0.162875), (61008,-0.189291), (61009,-0.326257), (61010,0.000798), (61011,0.241930), (61012,0.179277), (61013,0.020946), (61014,0.135731), (61015,0.047067), (61016,-0.077357), (61017,0.195823), (61018,0.070466), (61019,0.005490), (61020,0.271707), (61021,0.307995), (61022,0.168236), (61023,0.073073), (61024,-0.147042), (61025,0.151685), (61026,-0.012688), (61027,-0.018673), (61028,0.202948), (61029,0.327958), (61030,0.199808), (61031,0.140875), (61032,-0.003524), (61033,-0.156752), (61034,0.087631), (61035,0.348268), (61036,0.267037), (61037,0.122175), (61038,0.144061), (61039,-0.083486), (61040,-0.137773), (61041,-0.290068), (61042,-0.015035), (61043,0.208909), (61044,0.166701), (61045,0.004181), (61046,0.173780), (61047,0.140394), (61048,-0.100159), (61049,-0.259886), (61050,0.052773), (61051,0.266962), (61052,0.180621), (61053,0.017174), (61054,0.029775), (61055,-0.157823), (61056,-0.485702), (61057,-0.642179), (61058,0.055548), (61059,-0.065163), (61060,-0.112481), (61061,-0.299615), (61062,-0.047343), (61063,-0.176877), (61064,-0.350543), (61065,-0.380679), (61066,-0.123754), (61067,0.154072), (61068,-0.012625), (61069,-0.096179), (61070,-0.251730), (61071,-0.241453), (61072,-0.414186), (61073,-0.432249), (61074,-0.188793), (61075,0.120153), (61076,-0.041897), (61077,-0.103623), (61078,-0.195537), (61079,-0.032437), (61080,-0.156404), (61081,-0.211624), (61082,-0.368102), (61083,0.288286), (61084,0.134595), (61085,0.128153), (61086,-0.051086), (61087,-0.052424), (61088,-0.178244), (61089,-0.251116), (61090,-0.429885), (61091,0.249727), (61092,0.090463), (61093,0.039420), (61094,-0.088254), (61095,0.128721), (61096,-0.172213), (61097,-0.259950), (61098,0.019272), (61099,0.286409), (61100,0.122962), (61101,0.061242), (61102,-0.146330), (61103,-0.133730), (61104,-0.281385), (61105,-0.302228), (61106,-0.091753), (61107,0.186536), (61108,0.063032), (61109,-0.001937), (61110,-0.054834), (61111,0.094327), (61112,-0.324126), (61113,-0.374700), (61114,-0.147506), (61115,0.156794), (61116,0.018895), (61117,-0.105529), (61118,-0.287091), (61119,-0.276814), (61120,-0.430042), (61121,-0.473183), (61122,-0.198607), (61123,0.080145), (61124,-0.088411), (61125,-0.147344), (61126,-0.201631), (61127,-0.083597), (61128,-0.261903), (61129,-0.309227), (61130,-0.065771), (61131,0.202299), (61132,-0.006207), (61133,0.010576), (61134,-0.190960), (61135,-0.171397), (61136,-0.307900), (61137,-0.337109), (61138,-0.133133), (61139,0.147942), (61140,-0.016431), (61141,-0.068865), (61142,-0.157065), (61143,0.013930), (61144,-0.164382), (61145,-0.227961), (61146,-0.401627), (61147,0.276132), (61148,0.143806), (61149,0.093232), (61150,-0.086934), (61151,-0.068297), (61152,-0.222452), (61153,-0.281385), (61154,-0.384451), (61155,0.313277), (61156,0.129862), (61157,0.066746), (61158,-0.068831), (61159,0.129103), (61160,-0.012973), (61161,-0.070980), (61162,-0.211202), (61163,0.499068), (61164,0.332371), (61165,0.286443), (61166,0.116497), (61167,0.077532), (61168,-0.059897), (61169,-0.104898), (61170,-0.265559), (61171,0.396865), (61172,0.256186), (61173,0.233946), (61174,0.078395), (61175,0.269359), (61176,0.032989), (61177,-0.021298), (61178,-0.159197), (61179,0.530171), (61180,0.372297), (61181,0.312431), (61182,0.188470), (61183,0.160657), (61184,-0.034837), (61185,-0.083551), (61186,-0.234919), (61187,0.450267), (61188,0.306794), (61189,0.293847), (61190,0.122504), (61191,0.375246), (61192,0.081738), (61193,-0.022711), (61194,-0.176403), (61195,0.487881), (61196,0.303996), (61197,0.266891), (61198,0.101591), (61199,0.099789), (61200,-0.102211), (61201,-0.130023), (61202,-0.299970), (61203,0.370814), (61204,0.257535), (61205,0.185133), (61206,0.081141), (61207,0.286507), (61208,-0.049267), (61209,-0.220147), (61210,0.061399), (61211,0.303921), (61212,0.212934), (61213,0.042988), (61214,0.044436), (61215,-0.099499), (61216,-0.162152), (61217,-0.344177), (61218,-0.072851), (61219,0.178958), (61220,0.134426), (61221,0.012319), (61222,0.155907), (61223,0.101150), (61224,0.006914), (61225,-0.184861), (61226,0.079490), (61227,0.327122), (61228,0.275621), (61229,0.141442), (61230,0.139640), (61231,0.007777), (61232,-0.072521), (61233,-0.209957), (61234,0.033962), (61235,0.326184), (61236,0.251458), (61237,0.123315), (61238,0.267830), (61239,0.182879), (61240,0.031048), (61241,-0.143545), (61242,0.189553), (61243,0.367511), (61244,0.313224), (61245,0.163716), (61246,0.187462), (61247,-0.012678), (61248,-0.057679), (61249,-0.219266), (61250,0.058096), (61251,0.342885), (61252,0.280239), (61253,0.128401), (61254,0.288244), (61255,0.215379), (61256,0.057042), (61257,-0.079931), (61258,0.179780), (61259,0.368884), (61260,0.384271), (61261,0.228726), (61262,0.225065), (61263,0.048149), (61264,-0.014967), (61265,-0.187236), (61266,0.074328), (61267,0.333112), (61268,0.299257), (61269,0.101903), (61270,0.243168), (61271,0.177735), (61272,-0.037733), (61273,-0.193748), (61274,0.078962), (61275,0.289438), (61276,0.278350), (61277,0.126049), (61278,0.113565), (61279,-0.046163), (61280,-0.062830), (61281,-0.225343), (61282,0.019966), (61283,0.306151), (61284,0.243961), (61285,0.135793), (61286,0.244078), (61287,0.160523), (61288,0.018448), (61289,-0.085544), (61290,0.539723), (61291,0.386032), (61292,0.353109), (61293,0.179444), (61294,0.144668), (61295,-0.035504), (61296,-0.076322), (61297,-0.224434), (61298,0.417552), (61299,0.303341), (61300,0.243018), (61301,0.073998), (61302,0.344391), (61303,0.170725), (61304,-0.164122), (61305,-0.320130), (61306,0.343220), (61307,0.176524), (61308,0.149644), (61309,-0.009626), (61310,0.002511), (61311,-0.170222), (61312,0.117353), (61313,0.048664), (61314,0.267499), (61315,0.612675), (61316,0.414395), (61317,0.336877), (61318,0.254256), (61319,0.417349), (61320,0.050924), (61321,0.406783), (61322,0.262847), (61323,0.530448), (61324,0.400451), (61325,0.294599), (61326,0.106537), (61327,0.156758), (61328,-0.011799), (61329,0.343133), (61330,0.200594), (61331,0.438007), (61332,0.321010), (61333,0.324781), (61334,0.173876), (61335,0.284484), (61336,0.188394), (61337,0.110876), (61338,0.367801), (61339,0.637731), (61340,0.480320), (61341,0.456690), (61342,0.296956), (61343,0.282149), (61344,0.162835), (61345,0.101578), (61346,0.332022), (61347,0.601489), (61348,0.413421), (61349,0.372139), (61350,0.348510), (61351,0.466080), (61352,0.068998), (61353,0.371902), (61354,0.210315), (61355,0.509042), (61356,0.321444), (61357,0.246719), (61358,0.130185), (61359,0.146961), (61360,-0.025308), (61361,0.340306), (61362,0.162001), (61363,0.455149), (61364,0.303317), (61365,0.313131), (61366,0.167336), (61367,0.312314), (61368,0.158623), (61369,0.097830), (61370,0.304122), (61371,0.622361), (61372,0.507687), (61373,0.439461), (61374,0.238857), (61375,0.253781), (61376,0.116808), (61377,0.081563), (61378,0.259521), (61379,0.541993), (61380,0.372974), (61381,0.332156), (61382,0.263003), (61383,0.411695), (61384,0.049909), (61385,0.380690), (61386,0.209811), (61387,0.511324), (61388,0.357170), (61389,0.253641), (61390,0.045142), (61391,0.110690), (61392,0.025746), (61393,0.341199), (61394,0.165210), (61395,0.463010), (61396,0.351585), (61397,0.388337), (61398,0.292240), (61399,0.405171), (61400,0.237085), (61401,0.188364), (61402,0.422528), (61403,0.664587), (61404,0.547589), (61405,0.484479), (61406,0.294558), (61407,0.330846), (61408,0.194800), (61409,0.150732), (61410,0.333800), (61411,0.625558), (61412,0.456075), (61413,0.412007), (61414,0.378152), (61415,0.492010), (61416,0.434936), (61417,0.293787), (61418,0.626885), (61419,0.427678), (61420,0.704107), (61421,0.606621), (61422,0.466862), (61423,0.343365), (61424,0.355495), (61425,0.224102), (61426,0.528402), (61427,0.367748), (61428,0.649287), (61429,0.491877), (61430,0.520732), (61431,0.423246), (61432,0.373141), (61433,0.309562), (61434,0.579955), (61435,0.826654), (61436,0.657171), (61437,0.589415), (61438,0.401811), (61439,0.437172), (61440,0.284408), (61441,0.243127), (61442,0.506550), (61443,0.759292), (61444,0.597705), (61445,0.559210), (61446,0.494704), (61447,0.685668), (61448,0.488777), (61449,0.322544), (61450,0.688622), (61451,0.494055), (61452,0.769557), (61453,0.595898), (61454,0.537891), (61455,0.380950), (61456,0.374039), (61457,0.205020), (61458,0.598968), (61459,0.464319), (61460,0.700342), (61461,0.561509), (61462,0.624741), (61463,0.434357), (61464,0.238393), (61465,0.062411), (61466,0.755029), (61467,0.585076), (61468,0.543331), (61469,0.365952), (61470,0.383192), (61471,0.220678), (61472,0.153849), (61473,0.001085), (61474,0.679770), (61475,0.503781), (61476,0.481078), (61477,0.337143), (61478,0.561550), (61479,0.392531), (61480,0.318732), (61481,0.289993), (61482,0.519510), (61483,0.836352), (61484,0.662223), (61485,0.638587), (61486,0.470500), (61487,0.460802), (61488,0.300142), (61489,0.251891), (61490,0.502773), (61491,0.815902), (61492,0.633877), (61493,0.544287), (61494,0.516937), (61495,0.634045), (61496,0.331251), (61497,0.205894), (61498,0.918023), (61499,0.726705), (61500,0.662199), (61501,0.489466), (61502,0.476049), (61503,0.340943), (61504,0.315917), (61505,0.141324), (61506,0.821863), (61507,0.680251), (61508,0.581368), (61509,0.430000), (61510,0.696211), (61511,0.521155), (61512,0.397657), (61513,0.309920), (61514,0.555236), (61515,0.840488), (61516,0.690046), (61517,0.639479), (61518,0.477422), (61519,0.487236), (61520,0.321003), (61521,0.285294), (61522,0.530603), (61523,0.795887), (61524,0.622221), (61525,0.581403), (61526,0.523866), (61527,0.685563), (61528,0.318674), (61529,0.169160), (61530,0.839486), (61531,0.661637), (61532,0.614783), (61533,0.488493), (61534,0.429096), (61535,0.298630), (61536,0.233197), (61537,0.093901), (61538,0.773050), (61539,0.574300), (61540,0.524659), (61541,0.385370), (61542,0.682238), (61543,0.520651), (61544,0.218783), (61545,0.526339), (61546,0.388904), (61547,0.689491), (61548,0.531153), (61549,0.444349), (61550,0.324102), (61551,0.282820), (61552,0.096612), (61553,0.467800), (61554,0.308999), (61555,0.573820), (61556,0.442890), (61557,0.484287), (61558,0.341742), (61559,0.453740), (61560,0.276824), (61561,0.262480), (61562,0.478528), (61563,0.791658), (61564,0.658868), (61565,0.603185), (61566,0.413263), (61567,0.441656), (61568,0.219218), (61569,0.078532), (61570,0.606255), (61571,0.447454), (61572,0.403850), (61573,0.288712), (61574,0.635284), (61575,0.495062), (61576,0.351127), (61577,0.201612), (61578,0.599743), (61579,0.390311), (61580,0.301184), (61581,0.173974), (61582,0.398844), (61583,0.264195), (61584,0.210371), (61585,0.071545), (61586,0.614134), (61587,0.494813), (61588,0.415905), (61589,0.228770), (61590,0.598567), (61591,0.482966), (61592,0.300008), (61593,0.257800), (61594,0.487317), (61595,0.537074), (61596,0.405211), (61597,0.310511), (61598,0.136382), (61599,0.427676), (61600,0.255407), (61601,0.199723), (61602,0.432960), (61603,0.616028), (61604,0.423784), (61605,0.406190), (61606,0.344001), (61607,0.651557), (61608,0.193154), (61609,0.539263), (61610,0.369311), (61611,0.412568), (61612,0.231006), (61613,0.171146), (61614,-0.014135), (61615,0.267410), (61616,0.064947), (61617,0.393398), (61618,0.269901), (61619,0.425562), (61620,0.276517), (61621,0.324420), (61622,0.144249), (61623,0.414178), (61624,0.206606), (61625,0.176006), (61626,0.437107), (61627,0.497553), (61628,0.337356), (61629,0.312330), (61630,0.104294), (61631,0.382119), (61632,0.199161), (61633,0.137905), (61634,0.367892), (61635,0.522156), (61636,0.368934), (61637,0.328110), (61638,0.257104), (61639,0.547936), (61640,0.324101), (61641,0.315337), (61642,0.538811), (61643,0.550015), (61644,0.366136), (61645,0.273759), (61646,0.132141), (61647,0.404857), (61648,0.263708), (61649,0.226140), (61650,0.401312), (61651,0.570911), (61652,0.420933), (61653,0.362463), (61654,0.278445), (61655,0.581356), (61656,0.270202), (61657,0.197794), (61658,0.396190), (61659,0.440374), (61660,0.282507), (61661,0.262590), (61662,0.105180), (61663,0.358391), (61664,0.220028), (61665,0.168521), (61666,0.419409), (61667,0.566711), (61668,0.384222), (61669,0.357336), (61670,0.316518), (61671,0.572973), (61672,0.410459), (61673,0.349203), (61674,0.598225), (61675,0.562986), (61676,0.365632), (61677,0.398664), (61678,0.232431), (61679,0.500971), (61680,0.357029), (61681,0.290663), (61682,0.528546), (61683,0.651689), (61684,0.477097), (61685,0.450681), (61686,0.420545), (61687,0.701157), (61688,0.397900), (61689,0.348252), (61690,0.573587), (61691,0.599192), (61692,0.474768), (61693,0.400500), (61694,0.185501), (61695,0.448462), (61696,0.352829), (61697,0.236764), (61698,0.508084), (61699,0.647489), (61700,0.467787), (61701,0.387953), (61702,0.349921), (61703,0.635643), (61704,0.328202), (61705,0.267409), (61706,0.488104), (61707,0.539251), (61708,0.349793), (61709,0.310371), (61710,0.128346), (61711,0.402452), (61712,0.241329), (61713,0.181932), (61714,0.411449), (61715,0.553178), (61716,0.395304), (61717,0.383753), (61718,0.328069), (61719,0.615644), (61720,0.462886), (61721,0.307335), (61722,0.307393), (61723,0.510436), (61724,0.477514), (61725,0.302921), (61726,0.563559), (61727,0.416367), (61728,0.379732), (61729,0.234864), (61730,0.418395), (61731,0.612615), (61732,0.575047), (61733,0.382802), (61734,0.696395), (61735,0.682514), (61736,0.445681), (61737,0.269692), (61738,0.674323), (61739,0.561971), (61740,0.534159), (61741,0.358639), (61742,0.574687), (61743,0.460476), (61744,0.410829), (61745,0.221841), (61746,0.790903), (61747,0.654394), (61748,0.554122), (61749,0.367920), (61750,0.707987), (61751,0.634652), (61752,0.413147), (61753,0.282210), (61754,0.699853), (61755,0.560094), (61756,0.475613), (61757,0.315886), (61758,0.567231), (61759,0.385206), (61760,0.307695), (61761,0.139138), (61762,0.684049), (61763,0.535468), (61764,0.478858), (61765,0.312155), (61766,0.693098), (61767,0.576570), (61768,0.407087), (61769,0.213446), (61770,0.652917), (61771,0.503872), (61772,0.403600), (61773,0.306107), (61774,0.577896), (61775,0.406554), (61776,0.316500), (61777,0.157236), (61778,0.694245), (61779,0.540554), (61780,0.497413), (61781,0.367409), (61782,0.695867), (61783,0.534280), (61784,0.487889), (61785,0.327229), (61786,0.391387), (61787,0.645056), (61788,0.618639), (61789,0.436145), (61790,0.698178), (61791,0.510580), (61792,0.435855), (61793,0.286341), (61794,0.458726), (61795,0.688707), (61796,0.653461), (61797,0.521605), (61798,0.798497), (61799,0.723309), (61800,0.288137), (61801,0.541342), (61802,0.552546), (61803,0.421616), (61804,0.349207), (61805,0.163006), (61806,0.440362), (61807,0.304322), (61808,0.246322), (61809,0.459578), (61810,0.623141), (61811,0.420208), (61812,0.359884), (61813,0.283299), (61814,0.583880), (61815,0.388849), (61816,0.321557), (61817,0.180871), (61818,0.577606), (61819,0.417879), (61820,0.380311), (61821,0.245661), (61822,0.544858), (61823,0.365150), (61824,0.186381), (61825,0.118155), (61826,0.374616), (61827,0.555824), (61828,0.402133), (61829,0.335768), (61830,0.229916), (61831,0.486377), (61832,0.272298), (61833,0.191073), (61834,0.467503), (61835,0.460591), (61836,0.297145), (61837,0.281874), (61838,0.073838), (61839,0.376748), (61840,0.205869), (61841,0.200347), (61842,0.428938), (61843,0.582282), (61844,0.421621), (61845,0.388236), (61846,0.280061), (61847,0.536058), (61848,0.195174), (61849,0.172471), (61850,0.422890), (61851,0.428984), (61852,0.246496), (61853,0.236334), (61854,0.029688), (61855,0.295435), (61856,0.146854), (61857,0.112542), (61858,0.343918), (61859,0.494469), (61860,0.311981), (61861,0.276736), (61862,0.192718), (61863,0.472867), (61864,0.370735), (61865,0.197995), (61866,0.545031), (61867,0.427107), (61868,0.456889), (61869,0.273474), (61870,0.151367), (61871,-0.006971), (61872,0.323810), (61873,0.158040), (61874,0.513899), (61875,0.377396), (61876,0.523301), (61877,0.327807), (61878,0.416117), (61879,0.242458), (61880,0.340054), (61881,0.227239), (61882,0.561270), (61883,0.405255), (61884,0.444330), (61885,0.267878), (61886,0.232169), (61887,0.056180), (61888,0.318677), (61889,0.158950), (61890,0.503200), (61891,0.371800), (61892,0.515388), (61893,0.351478), (61894,0.324592), (61895,0.170901), (61896,0.439434), (61897,0.272274), (61898,0.609091), (61899,0.468406), (61900,0.426191), (61901,0.331961), (61902,0.213567), (61903,0.093319), (61904,0.370219), (61905,0.238825), (61906,0.594221), (61907,0.447029), (61908,0.580398), (61909,0.433207), (61910,0.467635), (61911,0.317200), (61912,0.353488), (61913,0.132910), (61914,0.454392), (61915,0.285372), (61916,0.321660), (61917,0.156824), (61918,0.087208), (61919,-0.025607), (61920,0.215519), (61921,0.049286), (61922,0.417224), (61923,0.248667), (61924,0.399688), (61925,0.274794), (61926,0.317588), (61927,0.171330), (61928,0.413383), (61929,0.274557), (61930,0.622983), (61931,0.473938), (61932,0.465637), (61933,0.278502), (61934,0.218636), (61935,0.076560), (61936,0.349740), (61937,0.218347), (61938,0.573742), (61939,0.387997), (61940,0.522756), (61941,0.395546), (61942,0.396994), (61943,0.247949), (61944,0.468174), (61945,0.283826), (61946,0.668025), (61947,0.526406), (61948,0.516245), (61949,0.362554), (61950,0.250202), (61951,0.114626), (61952,0.446797), (61953,0.322373), (61954,0.627137), (61955,0.464153), (61956,0.625393), (61957,0.500499), (61958,0.547470), (61959,0.356152), (61960,0.510423), (61961,0.355805), (61962,0.677757), (61963,0.542644), (61964,0.510185), (61965,0.331880), (61966,0.270623), (61967,0.122505), (61968,0.358991), (61969,0.213660), (61970,0.546294), (61971,0.403748), (61972,0.545013), (61973,0.408047), (61974,0.428537), (61975,0.277169), (61976,0.476029), (61977,0.447753), (61978,0.288952), (61979,0.661536), (61980,0.491120), (61981,0.429400), (61982,0.276642), (61983,0.530774), (61984,0.431428), (61985,0.392006), (61986,0.226236), (61987,0.771611), (61988,0.625352), (61989,0.528329), (61990,0.332835), (61991,0.754648), (61992,0.333408), (61993,0.287481), (61994,0.550441), (61995,0.571864), (61996,0.397741), (61997,0.362496), (61998,0.169319), (61999,0.440175), (62000,0.316678), (62001,0.254032), (62002,0.523028), (62003,0.654074), (62004,0.479482), (62005,0.435408), (62006,0.354177), (62007,0.637575), (62008,0.387736), (62009,0.325553), (62010,0.501652), (62011,0.548159), (62012,0.379603), (62013,0.319273), (62014,0.151186), (62015,0.428543), (62016,0.254413), (62017,0.200126), (62018,0.461697), (62019,0.610852), (62020,0.410711), (62021,0.384758), (62022,0.338831), (62023,0.623156), (62024,0.383073), (62025,0.308348), (62026,0.551334), (62027,0.536526), (62028,0.369366), (62029,0.317859), (62030,0.140017), (62031,0.435958), (62032,0.279944), (62033,0.236339), (62034,0.489544), (62035,0.630346), (62036,0.519384), (62037,0.464634), (62038,0.398268), (62039,0.665405), (62040,0.533085), (62041,0.493657), (62042,0.276798), (62043,0.698611), (62044,0.590443), (62045,0.518967), (62046,0.335552), (62047,0.613371), (62048,0.421127), (62049,0.422118), (62050,0.293042), (62051,0.791041), (62052,0.669397), (62053,0.642980), (62054,0.466065), (62055,0.854897), (62056,0.460138), (62057,0.397949), (62058,0.648837), (62059,0.610805), (62060,0.492411), (62061,0.425119), (62062,0.230551), (62063,0.554363), (62064,0.386740), (62065,0.305972), (62066,0.539202), (62067,0.701832), (62068,0.553720), (62069,0.446941), (62070,0.380112), (62071,0.659792), (62072,0.371863), (62073,0.346836), (62074,0.605614), (62075,0.640049), (62076,0.477992), (62077,0.391658), (62078,0.250972), (62079,0.508360), (62080,0.100589), (62081,-0.002940), (62082,0.287892), (62083,0.481642), (62084,0.251778), (62085,0.182625), (62086,0.166885), (62087,0.465612), (62088,0.280337), (62089,0.216295), (62090,0.444415), (62091,0.456552), (62092,0.294032), (62093,0.201192), (62094,0.062366), (62095,0.336472), (62096,0.139582), (62097,0.101550), (62098,0.342219), (62099,0.470473), (62100,0.345585), (62101,0.285256), (62102,0.240255), (62103,0.492996), (62104,0.211110), (62105,0.070424), (62106,0.418850), (62107,0.255867), (62108,0.296338), (62109,0.113380), (62110,0.038191), (62111,-0.108531), (62112,0.140491), (62113,0.007702), (62114,0.352415), (62115,0.222881), (62116,0.365536), (62117,0.193267), (62118,0.239304), (62119,0.089333), (62120,0.298875), (62121,0.149367), (62122,0.522877), (62123,0.325523), (62124,0.338587), (62125,0.216943), (62126,0.154760), (62127,0.002459), (62128,0.276572), (62129,0.117308), (62130,0.466661), (62131,0.315756), (62132,0.464454), (62133,0.323305), (62134,0.373062), (62135,0.200329), (62136,0.226398), (62137,0.092675), (62138,0.414164), (62139,0.286483), (62140,0.275396), (62141,0.157471), (62142,0.047906), (62143,-0.084883), (62144,0.179474), (62145,-0.004875), (62146,0.354697), (62147,0.226090), (62148,0.357600), (62149,0.177434), (62150,0.235087), (62151,0.098584), (62152,0.403348), (62153,0.253370), (62154,0.542811), (62155,0.419308), (62156,0.427725), (62157,0.303764), (62158,0.207205), (62159,0.050727), (62160,0.322517), (62161,0.134449), (62162,0.487521), (62163,0.332903), (62164,0.460700), (62165,0.317691), (62166,0.387886), (62167,0.197502), (62168,0.234253), (62169,0.101927), (62170,0.419232), (62171,0.249286), (62172,0.298579), (62173,0.068709), (62174,0.046932), (62175,-0.136483), (62176,0.144129), (62177,0.019236), (62178,0.355589), (62179,0.223263), (62180,0.338047), (62181,0.216410), (62182,0.244339), (62183,0.079959), (62184,0.348029), (62185,0.200380), (62186,0.520936), (62187,0.394189), (62188,0.386814), (62189,0.261457), (62190,0.151429), (62191,-0.067296), (62192,0.255589), (62193,0.126512), (62194,0.487017), (62195,0.341222), (62196,0.464835), (62197,0.301389), (62198,0.363224), (62199,0.222075), (62200,0.584903), (62201,0.438645), (62202,0.398290), (62203,0.569743), (62204,0.568874), (62205,0.459772), (62206,0.389693), (62207,0.238789), (62208,0.638773), (62209,0.486015), (62210,0.450300), (62211,0.657526), (62212,0.802041), (62213,0.620015), (62214,0.601958), (62215,0.469632), (62216,0.625756), (62217,0.445127), (62218,0.358787), (62219,0.602706), (62220,0.673364), (62221,0.491339), (62222,0.450521), (62223,0.261526), (62224,0.571406), (62225,0.377765), (62226,0.319758), (62227,0.562751), (62228,0.730490), (62229,0.560537), (62230,0.512750), (62231,0.493303), (62232,0.502647), (62233,0.415380), (62234,0.299315), (62235,0.674215), (62236,0.564187), (62237,0.494108), (62238,0.345057), (62239,0.617773), (62240,0.447363), (62241,0.386107), (62242,0.199436), (62243,0.779181), (62244,0.571608), (62245,0.547978), (62246,0.387781), (62247,0.754328), (62248,0.378141), (62249,0.331287), (62250,0.550585), (62251,0.544137), (62252,0.350503), (62253,0.305038), (62254,0.166206), (62255,0.451465), (62256,0.270836), (62257,0.204933), (62258,0.452102), (62259,0.618445), (62260,0.450358), (62261,0.394675), (62262,0.283250), (62263,0.564326), (62264,0.445011), (62265,0.383755), (62266,0.255142), (62267,0.673711), (62268,0.508874), (62269,0.457367), (62270,0.288818), (62271,0.542022), (62272,0.381825), (62273,0.349373), (62274,0.161305), (62275,0.715039), (62276,0.565531), (62277,0.530749), (62278,0.364516), (62279,0.762647), (62280,0.527667), (62281,0.451552), (62282,0.317366), (62283,0.667188), (62284,0.539508), (62285,0.485684), (62286,0.344535), (62287,0.603313), (62288,0.443122), (62289,0.389762), (62290,0.207737), (62291,0.736850), (62292,0.570153), (62293,0.523762), (62294,0.380290), (62295,0.764020), (62296,0.523003), (62297,0.432486), (62298,0.277399), (62299,0.719193), (62300,0.562715), (62301,0.495416), (62302,0.334762), (62303,0.607472), (62304,0.476079), (62305,0.385562), (62306,0.242553), (62307,0.801397), (62308,0.660248), (62309,0.593419), (62310,0.450873), (62311,0.802556), (62312,0.419399), (62313,0.334918), (62314,0.572331), (62315,0.635100), (62316,0.479086), (62317,0.418293), (62318,0.252986), (62319,0.546141), (62320,0.392450), (62321,0.319584), (62322,0.562107), (62323,0.681074), (62324,0.523664), (62325,0.467517), (62326,0.428558), (62327,0.730072), (62328,0.289321), (62329,0.223888), (62330,0.454332), (62331,0.450207), (62332,0.333679), (62333,0.293787), (62334,0.125694), (62335,0.355681), (62336,0.218245), (62337,0.121686), (62338,0.055783), (62339,0.580720), (62340,0.426565), (62341,0.395503), (62342,0.231593), (62343,0.612066), (62344,0.355727), (62345,0.295861), (62346,0.135671), (62347,0.539838), (62348,0.395433), (62349,0.321171), (62350,0.202320), (62351,0.396070), (62352,0.245629), (62353,0.209457), (62354,0.073881), (62355,0.582556), (62356,0.472064), (62357,0.372255), (62358,0.231106), (62359,0.622268), (62360,0.446749), (62361,0.299557), (62362,0.232728), (62363,0.495689), (62364,0.499923), (62365,0.291887), (62366,0.281726), (62367,0.116426), (62368,0.414220), (62369,0.233128), (62370,0.182554), (62371,0.396742), (62372,0.576091), (62373,0.375024), (62374,0.373686), (62375,0.303607), (62376,0.329676), (62377,0.173192), (62378,0.484925), (62379,0.300583), (62380,0.295061), (62381,0.111646), (62382,0.036451), (62383,-0.069858), (62384,0.187530), (62385,0.025473), (62386,0.396661), (62387,0.199777), (62388,0.366120), (62389,0.222648), (62390,0.198085), (62391,0.109427), (62392,0.342658), (62393,0.209868), (62394,0.130033), (62395,0.382312), (62396,0.399088), (62397,0.231002), (62398,0.177172), (62399,-0.013213), (62400,0.298520), (62401,0.111385), (62402,0.086822), (62403,0.374404), (62404,0.545856), (62405,0.361045), (62406,0.314190), (62407,0.247824), (62408,0.435075), (62409,0.263732), (62410,0.254961), (62411,0.490051), (62412,0.514730), (62413,0.352210), (62414,0.305819), (62415,0.160024), (62416,0.467574), (62417,0.265117), (62418,0.189922), (62419,0.406434), (62420,0.607617), (62421,0.422342), (62422,0.360622), (62423,0.284037), (62424,0.411364), (62425,0.257673), (62426,0.199666), (62427,0.478882), (62428,0.458039), (62429,0.303421), (62430,0.246811), (62431,0.034128), (62432,0.338892), (62433,0.201456), (62434,0.145773), (62435,0.392941), (62436,0.564864), (62437,0.413496), (62438,0.358275), (62439,0.323494), (62440,0.559980), (62441,0.413721), (62442,0.367794), (62443,0.598237), (62444,0.633135), (62445,0.519387), (62446,0.433053), (62447,0.233376), (62448,0.580876), (62449,0.403027), (62450,0.325979), (62451,0.576397), (62452,0.681432), (62453,0.517059), (62454,0.463699), (62455,0.416374), (62456,0.599906), (62457,0.418344), (62458,0.360344), (62459,0.607976), (62460,0.634045), (62461,0.455733), (62462,0.413055), (62463,0.234286), (62464,0.463333), (62465,0.330080), (62466,0.242813), (62467,0.484872), (62468,0.645642), (62469,0.502170), (62470,0.438127), (62471,0.317417), (62472,0.442890), (62473,0.304527), (62474,0.240015), (62475,0.507158), (62476,0.485382), (62477,0.341446), (62478,0.328962), (62479,0.179454), (62480,0.451701), (62481,0.241811), (62482,0.199133), (62483,0.428650), (62484,0.582451), (62485,0.410645), (62486,0.374473), (62487,0.327618), (62488,0.406636), (62489,0.341197), (62490,0.146166), (62491,0.584247), (62492,0.429160), (62493,0.355825), (62494,0.247193), (62495,0.469277), (62496,0.323018), (62497,0.230178), (62498,0.099242), (62499,0.641367), (62500,0.495108), (62501,0.428743), (62502,0.339152), (62503,0.701517), (62504,0.495334), (62505,0.427109), (62506,0.289679), (62507,0.659933), (62508,0.566167), (62509,0.503514), (62510,0.391162), (62511,0.612783), (62512,0.444697), (62513,0.363929), (62514,0.257150), (62515,0.744930), (62516,0.579160), (62517,0.551348), (62518,0.382328), (62519,0.753979), (62520,0.446545), (62521,0.363917), (62522,0.237170), (62523,0.615327), (62524,0.450484), (62525,0.371576), (62526,0.248542), (62527,0.482242), (62528,0.311362), (62529,0.258935), (62530,0.100598), (62531,0.632034), (62532,0.459764), (62533,0.443567), (62534,0.271298), (62535,0.645735), (62536,0.423297), (62537,0.342999), (62538,0.206490), (62539,0.596262), (62540,0.432351), (62541,0.391070), (62542,0.239232), (62543,0.519381), (62544,0.387525), (62545,0.299324), (62546,0.184186), (62547,0.729561), (62548,0.566114), (62549,0.461659), (62550,0.292639), (62551,0.711208), (62552,0.429779), (62553,0.323933), (62554,0.206936), (62555,0.627828), (62556,0.467168), (62557,0.377578), (62558,0.173718), (62559,0.449221), (62560,0.350344), (62561,0.231487), (62562,0.088948), (62563,0.656151), (62564,0.514069), (62565,0.444916), (62566,0.279153), (62567,0.685637), (62568,0.282049), (62569,0.233798), (62570,0.476321), (62571,0.482421), (62572,0.308755), (62573,0.239603), (62574,0.108673), (62575,0.355372), (62576,0.213297), (62577,0.191057), (62578,0.432183), (62579,0.591100), (62580,0.426263), (62581,0.377549), (62582,0.286098), (62583,0.584362), (62584,0.416269), (62585,0.343398), (62586,0.161842), (62587,0.560900), (62588,0.390484), (62589,0.322259), (62590,0.175074), (62591,0.475191), (62592,0.163574), (62593,0.113464), (62594,-0.025826), (62595,0.495861), (62596,0.372827), (62597,0.324576), (62598,0.182958), (62599,0.509556), (62600,0.387918), (62601,0.182199), (62602,0.086109), (62603,0.370434), (62604,0.391857), (62605,0.262787), (62606,0.208030), (62607,0.022755), (62608,0.326592), (62609,0.163609), (62610,0.094920), (62611,0.348131), (62612,0.447123), (62613,0.314334), (62614,0.256327), (62615,0.142586), (62616,0.318684), (62617,0.170103), (62618,0.128821), (62619,0.389922), (62620,0.390443), (62621,0.256727), (62622,0.188502), (62623,-0.010706), (62624,0.311710), (62625,0.188676), (62626,0.113018), (62627,0.339748), (62628,0.505164), (62629,0.355656), (62630,0.287894), (62631,0.247076), (62632,0.256889), (62633,0.104588), (62634,0.484605), (62635,0.296074), (62636,0.306351), (62637,0.120143), (62638,0.051924), (62639,-0.097591), (62640,0.232257), (62641,0.058597), (62642,0.360111), (62643,0.234754), (62644,0.367653), (62645,0.203280), (62646,0.244677), (62647,0.107705), (62648,0.390177), (62649,0.184927), (62650,0.129244), (62651,0.390814), (62652,0.404341), (62653,0.266905), (62654,0.168956), (62655,-0.013069), (62656,0.250818), (62657,0.139863), (62658,0.043766), (62659,0.288612), (62660,0.499087), (62661,0.344000), (62662,0.266488), (62663,0.181074), (62664,0.452864), (62665,0.267119), (62666,0.228161), (62667,0.454892), (62668,0.454017), (62669,0.313337), (62670,0.263690), (62671,0.109999), (62672,0.377606), (62673,0.199294), (62674,0.092985), (62675,0.370341), (62676,0.545050), (62677,0.412260), (62678,0.377948), (62679,0.260950), (62680,0.369235), (62681,0.200215), (62682,0.161720), (62683,0.397273), (62684,0.432635), (62685,0.299382), (62686,0.260417), (62687,0.069569), (62688,0.339499), (62689,0.229001), (62690,0.137557), (62691,0.361031), (62692,0.512052), (62693,0.300760), (62694,0.278057), (62695,0.252567), (62696,0.487194), (62697,0.340008), (62698,0.230907), (62699,0.498050), (62700,0.534338), (62701,0.404335), (62702,0.321714), (62703,0.097879), (62704,0.373382), (62705,0.211795), (62706,0.182123), (62707,0.468778), (62708,0.617005), (62709,0.438700), (62710,0.416460), (62711,0.364953), (62712,0.509938), (62713,0.352064), (62714,0.274552), (62715,0.550982), (62716,0.575654), (62717,0.377837), (62718,0.296606), (62719,0.109471), (62720,0.441179), (62721,0.276805), (62722,0.268967), (62723,0.514740), (62724,0.645322), (62725,0.478156), (62726,0.408540), (62727,0.353790), (62728,0.460215), (62729,0.294909), (62730,0.239225), (62731,0.482217), (62732,0.487379), (62733,0.346230), (62734,0.337465), (62735,0.149397), (62736,0.412358), (62737,0.249844), (62738,0.192771), (62739,0.426928), (62740,0.581198), (62741,0.430763), (62742,0.348136), (62743,0.307317), (62744,0.473667), (62745,0.424946), (62746,0.298199), (62747,0.301507), (62748,0.553785), (62749,0.511107), (62750,0.366709), (62751,0.644065), (62752,0.462040), (62753,0.418435), (62754,0.262884), (62755,0.436666), (62756,0.668969), (62757,0.619322), (62758,0.432188), (62759,0.726275), (62760,0.487575), (62761,0.406351), (62762,0.251263), (62763,0.667510), (62764,0.512885), (62765,0.387535), (62766,0.240807), (62767,0.558582), (62768,0.399781), (62769,0.313904), (62770,0.172755), (62771,0.713484), (62772,0.542141), (62773,0.509219), (62774,0.319297), (62775,0.719282), (62776,0.364003), (62777,0.297174), (62778,0.159738), (62779,0.579234), (62780,0.435299), (62781,0.364750), (62782,0.211522), (62783,0.466587), (62784,0.292458), (62785,0.264645), (62786,0.129539), (62787,0.663298), (62788,0.475236), (62789,0.402828), (62790,0.250070), (62791,0.628690), (62792,0.400679), (62793,0.341746), (62794,0.148569), (62795,0.553200), (62796,0.398118), (62797,0.326180), (62798,0.158087), (62799,0.413615), (62800,0.294764), (62801,0.218179), (62802,0.055659), (62803,0.592674), (62804,0.433873), (62805,0.423249), (62806,0.252833), (62807,0.667219), (62808,0.540003), (62809,0.499654), (62810,0.301367), (62811,0.345088), (62812,0.596903), (62813,0.524495), (62814,0.354085), (62815,0.642593), (62816,0.468001), (62817,0.397452), (62818,0.236792), (62819,0.417073), (62820,0.664242), (62821,0.601595), (62822,0.411674), (62823,0.703432), (62824,0.442441), (62825,0.278068), (62826,0.606056), (62827,0.412421), (62828,0.457069), (62829,0.324279), (62830,0.241188), (62831,0.084711), (62832,0.374615), (62833,0.210242), (62834,0.547059), (62835,0.402191), (62836,0.506293), (62837,0.342846), (62838,0.390286), (62839,0.282581), (62840,0.382963), (62841,0.319390), (62842,0.188923), (62843,0.561501), (62844,0.421279), (62845,0.413904), (62846,0.269969), (62847,0.466975), (62848,0.388530), (62849,0.220901), (62850,0.131310), (62851,0.447226), (62852,0.572230), (62853,0.410179), (62854,0.343350), (62855,0.234718), (62856,0.440541), (62857,0.258052), (62858,0.194009), (62859,0.459293), (62860,0.513233), (62861,0.319592), (62862,0.312681), (62863,0.143661), (62864,0.404305), (62865,0.268259), (62866,0.191675), (62867,0.473220), (62868,0.611692), (62869,0.444996), (62870,0.426475), (62871,0.343384), (62872,0.519953), (62873,0.326312), (62874,0.296176), (62875,0.538236), (62876,0.578706), (62877,0.381816), (62878,0.282470), (62879,0.130175), (62880,0.408928), (62881,0.242231), (62882,0.199090), (62883,0.449972), (62884,0.576835), (62885,0.452874), (62886,0.371643), (62887,0.262541), (62888,-0.025851), (62889,0.245006), (62890,0.524691), (62891,0.476441), (62892,0.323676), (62893,0.357641), (62894,0.144959), (62895,0.127365), (62896,-0.017967), (62897,0.274725), (62898,0.489376), (62899,0.434163), (62900,0.296727), (62901,0.467716), (62902,0.373479), (62903,0.317333), (62904,0.455811), (62905,0.273786), (62906,0.252010), (62907,0.544237), (62908,0.537789), (62909,0.325570), (62910,0.275460), (62911,0.096228), (62912,0.357328), (62913,0.179480), (62914,0.144241), (62915,0.424847), (62916,0.549856), (62917,0.411494), (62918,0.369279), (62919,0.299200), (62920,0.197068), (62921,0.450736), (62922,0.348604), (62923,0.706322), (62924,0.504322), (62925,0.457468), (62926,0.307490), (62927,0.208614), (62928,0.078610), (62929,0.331352), (62930,0.200422), (62931,0.550245), (62932,0.414668), (62933,0.556860), (62934,0.395736), (62935,0.428305), (62936,0.467849), (62937,0.314158), (62938,0.248719), (62939,0.505643), (62940,0.474575), (62941,0.354797), (62942,0.313046), (62943,0.085498), (62944,0.395377), (62945,0.262124), (62946,0.209227), (62947,0.410410), (62948,0.565144), (62949,0.371040), (62950,0.333472), (62951,0.263856), (62952,0.182625), (62953,0.453019), (62954,0.279353), (62955,0.633358), (62956,0.493136), (62957,0.494121), (62958,0.380842), (62959,0.364639), (62960,0.183547), (62961,0.441861), (62962,0.251013), (62963,0.621267), (62964,0.497307), (62965,0.654827), (62966,0.482094), (62967,0.517913), (62968,0.582071), (62969,0.430240), (62970,0.369447), (62971,0.572020), (62972,0.610168), (62973,0.454617), (62974,0.391507), (62975,0.196940), (62976,0.498917), (62977,0.357768), (62978,0.324383), (62979,0.561796), (62980,0.725352), (62981,0.516853), (62982,0.486254), (62983,0.416632), (62984,0.213242), (62985,0.459484), (62986,0.351778), (62987,0.697418), (62988,0.468011), (62989,0.488507), (62990,0.374765), (62991,0.258694), (62992,0.166317), (62993,0.406517), (62994,0.233784), (62995,0.590570), (62996,0.446171), (62997,0.579077), (62998,0.430495), (62999,0.449595), (63000,0.492846), (63001,0.344734), (63002,0.286727), (63003,0.566407), (63004,0.605018), (63005,0.393732), (63006,0.371955), (63007,0.149054), (63008,0.441745), (63009,0.286194), (63010,0.296935), (63011,0.532488), (63012,0.646345), (63013,0.479186), (63014,0.433721), (63015,0.417524), (63016,0.670265), (63017,0.518434), (63018,0.458105), (63019,0.677866), (63020,0.707185), (63021,0.586937), (63022,0.547515), (63023,0.340406), (63024,0.649352), (63025,0.496124), (63026,0.473421), (63027,0.684823), (63028,0.841880), (63029,0.697482), (63030,0.653407), (63031,0.544312), (63032,0.628902), (63033,0.451523), (63034,0.415351), (63035,0.640222), (63036,0.609160), (63037,0.471261), (63038,0.414650), (63039,0.283721), (63040,0.552717), (63041,0.360937), (63042,0.329874), (63043,0.521301), (63044,0.710405), (63045,0.527454), (63046,0.466197), (63047,0.364528), (63048,0.579186), (63049,0.401801), (63050,0.338222), (63051,0.580744), (63052,0.600777), (63053,0.435477), (63054,0.365855), (63055,0.147600), (63056,0.419389), (63057,0.277307), (63058,0.207228), (63059,0.492017), (63060,0.672298), (63061,0.522327), (63062,0.463857), (63063,0.358005), (63064,0.586132), (63065,0.465421), (63066,0.385117), (63067,0.629962), (63068,0.598900), (63069,0.473080), (63070,0.436901), (63071,0.240480), (63072,0.502045), (63073,0.335811), (63074,0.309395), (63075,0.537516), (63076,0.695969), (63077,0.532986), (63078,0.473126), (63079,0.386322), (63080,0.479278), (63081,0.342306), (63082,0.667977), (63083,0.514749), (63084,0.511551), (63085,0.356933), (63086,0.280812), (63087,0.137340), (63088,0.417489), (63089,0.251255), (63090,0.569024), (63091,0.388859), (63092,0.537093), (63093,0.421022), (63094,0.443378), (63095,0.270639), (63096,0.566580), (63097,0.419858), (63098,0.384613), (63099,0.572327), (63100,0.546837), (63101,0.421480), (63102,0.392734), (63103,0.220465), (63104,0.343615), (63105,0.144401), (63106,0.097077), (63107,0.354002), (63108,0.508736), (63109,0.383379), (63110,0.306330), (63111,0.249720), (63112,0.396088), (63113,0.269805), (63114,0.236419), (63115,0.476155), (63116,0.450202), (63117,0.309053), (63118,0.310965), (63119,0.132659), (63120,0.386327), (63121,0.230313), (63122,0.181599), (63123,0.441310), (63124,0.595111), (63125,0.383361), (63126,0.337434), (63127,0.249233), (63128,0.100188), (63129,0.402166), (63130,0.244761), (63131,0.571823), (63132,0.393511), (63133,0.437231), (63134,0.304905), (63135,0.224607), (63136,0.057910), (63137,0.325517), (63138,0.154638), (63139,0.510497), (63140,0.420906), (63141,0.555202), (63142,0.353665), (63143,0.413648), (63144,-0.018744), (63145,0.269764), (63146,0.483952), (63147,0.456603), (63148,0.309881), (63149,0.321085), (63150,0.132097), (63151,0.071767), (63152,-0.082387), (63153,0.205651), (63154,0.445857), (63155,0.389710), (63156,0.197930), (63157,0.356377), (63158,0.294657), (63159,0.216212), (63160,0.029078), (63161,0.309690), (63162,0.169937), (63163,0.509535), (63164,0.381861), (63165,0.382382), (63166,0.237977), (63167,0.133521), (63168,0.003055), (63169,0.274845), (63170,0.124403), (63171,0.411052), (63172,0.322858), (63173,0.481305), (63174,0.291847), (63175,0.325349), (63176,0.133104), (63177,0.427655), (63178,0.283713), (63179,0.617281), (63180,0.476595), (63181,0.467361), (63182,0.335034), (63183,0.242658), (63184,0.096863), (63185,0.378871), (63186,0.201492), (63187,0.521121), (63188,0.386472), (63189,0.516121), (63190,0.362900), (63191,0.423339), (63192,0.107540), (63193,0.345879), (63194,0.229815), (63195,0.584283), (63196,0.409684), (63197,0.426931), (63198,0.311329), (63199,0.208734), (63200,0.081980), (63201,0.350050), (63202,0.164312), (63203,0.459783), (63204,0.351614), (63205,0.537469), (63206,0.428837), (63207,0.461405), (63208,0.300282), (63209,0.540018), (63210,0.354279), (63211,0.689237), (63212,0.555984), (63213,0.558828), (63214,0.472488), (63215,0.375001), (63216,0.193903), (63217,0.493563), (63218,0.294813), (63219,0.620478), (63220,0.475616), (63221,0.625240), (63222,0.472012), (63223,0.533385), (63224,0.249632), (63225,0.536281), (63226,0.354256), (63227,0.676677), (63228,0.547601), (63229,0.575530), (63230,0.410223), (63231,0.288585), (63232,0.207354), (63233,0.440121), (63234,0.259956), (63235,0.596310), (63236,0.416138), (63237,0.604315), (63238,0.467349), (63239,0.502704), (63240,0.177155), (63241,0.499570), (63242,0.321258), (63243,0.691056), (63244,0.485336), (63245,0.523484), (63246,0.373043), (63247,0.301104), (63248,0.149736), (63249,0.377863), (63250,0.272474), (63251,0.581421), (63252,0.437485), (63253,0.575031), (63254,0.449674), (63255,0.435336), (63256,0.689468), (63257,0.528814), (63258,0.475917), (63259,0.324086), (63260,0.764014), (63261,0.597317), (63262,0.538384), (63263,0.353572), (63264,0.634648), (63265,0.470738), (63266,0.380221), (63267,0.221420), (63268,0.757039), (63269,0.604274), (63270,0.573675), (63271,0.413485), (63272,0.581224), (63273,0.436819), (63274,0.448023), (63275,0.662681), (63276,0.661342), (63277,0.525303), (63278,0.508636), (63279,0.303850), (63280,0.562634), (63281,0.419625), (63282,0.327248), (63283,0.593459), (63284,0.741687), (63285,0.588929), (63286,0.488186), (63287,0.427863), (63288,0.508277), (63289,0.370378), (63290,0.272892), (63291,0.560467), (63292,0.563781), (63293,0.410090), (63294,0.375771), (63295,0.203502), (63296,0.502692), (63297,0.333673), (63298,0.254765), (63299,0.515866), (63300,0.632516), (63301,0.475105), (63302,0.432891), (63303,0.324722), (63304,0.504540), (63305,0.375000), (63306,0.306312), (63307,0.576241), (63308,0.588842), (63309,0.455125), (63310,0.379004), (63311,0.221130), (63312,0.457616), (63313,0.307175), (63314,0.233840), (63315,0.466150), (63316,0.651534), (63317,0.501099), (63318,0.469104), (63319,0.359075), (63320,0.666162), (63321,0.549170), (63322,0.473049), (63323,0.296133), (63324,0.692405), (63325,0.539177), (63326,0.498822), (63327,0.315401), (63328,0.580221), (63329,0.442785), (63330,0.366200), (63331,0.232947), (63332,0.772286), (63333,0.611625), (63334,0.574990), (63335,0.402251), (63336,0.432966), (63337,0.269519), (63338,0.649536), (63339,0.474943), (63340,0.482427), (63341,0.328743), (63342,0.302320), (63343,0.147702), (63344,0.405553), (63345,0.300171), (63346,0.637915), (63347,0.485150), (63348,0.631525), (63349,0.455536), (63350,0.470923), (63351,0.325591), (63352,0.569510), (63353,0.421855), (63354,0.378714), (63355,0.625882), (63356,0.604106), (63357,0.438342), (63358,0.346892), (63359,0.231754), (63360,0.403207), (63361,0.299221), (63362,0.185473), (63363,0.409417), (63364,0.526524), (63365,0.355188), (63366,0.296718), (63367,0.226170), (63368,0.459869), (63369,0.320574), (63370,0.241203), (63371,0.481872), (63372,0.526982), (63373,0.355176), (63374,0.266049), (63375,0.097956), (63376,0.402256), (63377,0.220701), (63378,0.116245), (63379,0.356908), (63380,0.512105), (63381,0.353774), (63382,0.290195), (63383,0.214537), (63384,0.405037), (63385,0.263425), (63386,0.192413), (63387,0.440509), (63388,0.447530), (63389,0.267364), (63390,0.246521), (63391,0.089110), (63392,0.353004), (63393,0.201172), (63394,0.185432), (63395,0.360604), (63396,0.536239), (63397,0.396487), (63398,0.359382), (63399,0.279084), (63400,0.143971), (63401,0.457564), (63402,0.307586), (63403,0.642543), (63404,0.467950), (63405,0.460112), (63406,0.337079), (63407,0.233086), (63408,0.097510), (63409,0.327954), (63410,0.206316), (63411,0.570998), (63412,0.392229), (63413,0.546963), (63414,0.413710), (63415,0.439309), (63416,0.149990), (63417,0.433389), (63418,0.279698), (63419,0.624411), (63420,0.467463), (63421,0.440584), (63422,0.285960), (63423,0.203339), (63424,0.064049), (63425,0.316321), (63426,0.141729), (63427,0.543573), (63428,0.394065), (63429,0.524648), (63430,0.392785), (63431,0.415604), (63432,0.231256), (63433,0.475168), (63434,0.319624), (63435,0.631356), (63436,0.520395), (63437,0.546927), (63438,0.379304), (63439,0.287854), (63440,0.155534), (63441,0.412922), (63442,0.260621), (63443,0.607193), (63444,0.435851), (63445,0.559464), (63446,0.411809), (63447,0.475968), (63448,0.042649), (63449,0.300500), (63450,0.170960), (63451,0.529612), (63452,0.379634), (63453,0.363437), (63454,0.213459), (63455,0.133161), (63456,-0.013567), (63457,0.260545), (63458,0.057149), (63459,0.386070), (63460,0.221697), (63461,0.417770), (63462,0.268262), (63463,0.308263), (63464,0.146676), (63465,0.429611), (63466,0.279170), (63467,0.668936), (63468,0.478088), (63469,0.494401), (63470,0.296584), (63471,0.238114), (63472,0.125299), (63473,0.359463), (63474,0.189510), (63475,0.549551), (63476,0.404226), (63477,0.543625), (63478,0.382971), (63479,0.429941), (63480,0.401665), (63481,0.653474), (63482,0.513721), (63483,0.469184), (63484,0.675939), (63485,0.683430), (63486,0.545068), (63487,0.468019), (63488,0.460181), (63489,0.345507), (63490,0.233155), (63491,0.110585), (63492,0.648990), (63493,0.518523), (63494,0.415001), (63495,0.274315), (63496,0.143385), (63497,0.404023), (63498,0.235930), (63499,0.172351), (63500,0.418129), (63501,0.466490), (63502,0.285861), (63503,0.248293), (63504,0.076486), (63505,0.383573), (63506,0.232668), (63507,0.210429), (63508,0.418581), (63509,0.567278), (63510,0.427983), (63511,0.328173), (63512,0.445287), (63513,0.319467), (63514,0.263783), (63515,0.099410), (63516,0.511937), (63517,0.398189), (63518,0.295593), (63519,0.174419), (63520,0.448062), (63521,0.320845), (63522,0.252156), (63523,0.070131), (63524,0.605750), (63525,0.439053), (63526,0.415887), (63527,0.256160), (63528,0.317062), (63529,0.220972), (63530,0.118376), (63531,0.368795), (63532,0.392541), (63533,0.225844), (63534,0.191062), (63535,0.001604), (63536,0.285003), (63537,0.091369), (63538,0.040332), (63539,0.267062), (63540,0.484501), (63541,0.316408), (63542,0.270480), (63543,0.155805), (63544,0.481477), (63545,0.337071), (63546,0.247481), (63547,0.094260), (63548,0.476129), (63549,0.372137), (63550,0.338288), (63551,0.195743), (63552,0.459167), (63553,0.277611), (63554,0.251189), (63555,0.079846), (63556,0.578308), (63557,0.406039), (63558,0.365684), (63559,0.244503), (63560,0.540444), (63561,0.399759), (63562,0.339899), (63563,0.186671), (63564,0.633105), (63565,0.501712), (63566,0.367995), (63567,0.264466), (63568,0.467972), (63569,0.313818), (63570,0.234910), (63571,0.090511), (63572,0.645172), (63573,0.479408), (63574,0.471564), (63575,0.300228), (63576,0.561328), (63577,0.409027), (63578,0.382611), (63579,0.216841), (63580,0.599644), (63581,0.437124), (63582,0.413494), (63583,0.213817), (63584,0.488857), (63585,0.364896), (63586,0.243252), (63587,0.096530), (63588,0.631686), (63589,0.531876), (63590,0.439030), (63591,0.311350), (63592,0.462834), (63593,0.335154), (63594,0.279007), (63595,0.495055), (63596,0.520661), (63597,0.357214), (63598,0.289921), (63599,0.078166), (63600,0.394545), (63601,0.239457), (63602,0.207931), (63603,0.446271), (63604,0.613084), (63605,0.441741), (63606,0.377698), (63607,0.309009), (63608,0.468389), (63609,0.310979), (63610,0.216749), (63611,0.475063), (63612,0.439354), (63613,0.261969), (63614,0.223474), (63615,0.049345), (63616,0.026642), (63617,-0.128439), (63618,0.239961), (63619,0.082551), (63620,0.172721), (63621,-0.017664), (63622,0.063677), (63623,-0.103483), (63624,0.078658), (63625,-0.094081), (63626,0.244133), (63627,0.113203), (63628,0.146698), (63629,0.018554), (63630,-0.068713), (63631,-0.216361), (63632,0.063318), (63633,-0.087123), (63634,0.232975), (63635,0.064882), (63636,0.202891), (63637,0.062212), (63638,0.093854), (63639,-0.039399), (63640,-0.034702), (63641,0.221296), (63642,0.075031), (63643,0.391874), (63644,0.217281), (63645,0.218272), (63646,0.080373), (63647,0.014934), (63648,-0.140147), (63649,0.149751), (63650,-0.048993), (63651,0.301287), (63652,0.163394), (63653,0.320444), (63654,0.176509), (63655,0.187713), (63656,-0.134123), (63657,0.148349), (63658,0.402481), (63659,0.342621), (63660,0.184284), (63661,0.175049), (63662,0.019968), (63663,-0.075665), (63664,-0.207058), (63665,0.141831), (63666,0.331869), (63667,0.297556), (63668,0.054680), (63669,0.232175), (63670,0.163486), (63671,0.138923), (63672,-0.279993), (63673,-0.022142), (63674,0.236636), (63675,0.178635), (63676,-0.015469), (63677,0.025929), (63678,-0.169102), (63679,-0.243833), (63680,-0.387768), (63681,-0.069993), (63682,0.140939), (63683,0.100584), (63684,-0.104665), (63685,0.095591), (63686,0.007397), (63687,-0.009270), (63688,-0.272584), (63689,0.049831), (63690,0.316048), (63691,0.268260), (63692,0.095058), (63693,0.090939), (63694,-0.083190), (63695,-0.118435), (63696,-0.293961), (63697,-0.011489), (63698,0.240789), (63699,0.214367), (63700,0.036061), (63701,0.198691), (63702,0.121643), (63703,0.065496), (63704,-0.094701), (63705,0.189624), (63706,0.019678), (63707,0.303540), (63708,0.174470), (63709,0.206112), (63710,0.067749), (63711,0.000920), (63712,-0.171356), (63713,0.105080), (63714,-0.035142), (63715,0.273341), (63716,0.077840), (63717,0.227465), (63718,0.095145), (63719,0.088234), (63720,-0.050129), (63721,0.235130), (63722,0.119059), (63723,0.485136), (63724,0.335165), (63725,0.322217), (63726,0.151801), (63727,0.057101), (63728,-0.068719), (63729,0.219789), (63730,0.090249), (63731,0.335095), (63732,0.275235), (63733,0.415567), (63734,0.215427), (63735,0.256361), (63736,0.047392), (63737,0.329401), (63738,0.202184), (63739,0.553866), (63740,0.466592), (63741,0.470370), (63742,0.280449), (63743,0.172274), (63744,-0.031116), (63745,0.269934), (63746,0.095805), (63747,0.469315), (63748,0.301222), (63749,0.450847), (63750,0.283687), (63751,0.296750), (63752,-0.009757), (63753,0.255990), (63754,0.123201), (63755,0.450725), (63756,0.332338), (63757,0.338432), (63758,0.174522), (63759,0.090041), (63760,-0.024634), (63761,0.257375), (63762,0.086032), (63763,0.406124), (63764,0.263115), (63765,0.375583), (63766,0.264158), (63767,0.253997), (63768,0.235940), (63769,0.088749), (63770,0.049327), (63771,0.307178), (63772,0.332777), (63773,0.147039), (63774,0.099715), (63775,-0.121327), (63776,0.222460), (63777,0.041361), (63778,0.007043), (63779,0.221237), (63780,0.384330), (63781,0.188836), (63782,0.097850), (63783,0.011973), (63784,0.284225), (63785,0.143540), (63786,0.088790), (63787,0.337812), (63788,0.369453), (63789,0.234341), (63790,0.187486), (63791,-0.013581), (63792,0.246124), (63793,0.110084), (63794,0.022817), (63795,0.235616), (63796,0.408928), (63797,0.209714), (63798,0.229747), (63799,0.167558), (63800,0.339017), (63801,0.164424), (63802,0.120819), (63803,0.348477), (63804,0.369436), (63805,0.197630), (63806,0.141014), (63807,-0.003385), (63808,0.263295), (63809,0.097525), (63810,0.041378), (63811,0.282041), (63812,0.427019), (63813,0.280297), (63814,0.208822), (63815,0.161035), (63816,0.363151), (63817,0.189021), (63818,0.116150), (63819,0.363782), (63820,0.415398), (63821,0.245452), (63822,0.225072), (63823,-0.051248), (63824,0.298575), (63825,0.097038), (63826,0.089664), (63827,0.297353), (63828,0.472524), (63829,0.287713), (63830,0.283125), (63831,0.181456), (63832,0.292527), (63833,0.108179), (63834,0.037630), (63835,0.338680), (63836,0.349884), (63837,0.235679), (63838,0.138656), (63839,-0.034546), (63840,0.260468), (63841,0.124892), (63842,0.080354), (63843,0.316377), (63844,0.412583), (63845,0.253319), (63846,0.215751), (63847,0.191651), (63848,0.292040), (63849,0.180152), (63850,0.548089), (63851,0.347022), (63852,0.306668), (63853,0.162732), (63854,0.097756), (63855,-0.050362), (63856,0.218641), (63857,0.092821), (63858,0.413376), (63859,0.248540), (63860,0.404200), (63861,0.229608), (63862,0.234775), (63863,0.115918), (63864,0.118299), (63865,0.040787), (63866,0.386890), (63867,0.219267), (63868,0.203527), (63869,0.036367), (63870,-0.038822), (63871,-0.171611), (63872,-0.048468), (63873,-0.184037), (63874,0.158816), (63875,0.039495), (63876,0.121306), (63877,-0.036568), (63878,-0.006317), (63879,-0.168837), (63880,-0.022925), (63881,-0.168721), (63882,0.211753), (63883,0.052489), (63884,0.052084), (63885,-0.104394), (63886,-0.187948), (63887,-0.334207), (63888,-0.120018), (63889,-0.254661), (63890,0.059395), (63891,-0.072005), (63892,0.110136), (63893,-0.006861), (63894,-0.033747), (63895,-0.170714), (63896,0.152165), (63897,0.010089), (63898,-0.045131), (63899,0.232695), (63900,0.265733), (63901,0.087885), (63902,0.016409), (63903,-0.136818), (63904,0.163769), (63905,0.003108), (63906,-0.090195), (63907,0.166729), (63908,0.297305), (63909,0.157083), (63910,0.124161), (63911,-0.004446), (63912,-0.212482), (63913,0.041656), (63914,0.221468), (63915,0.210843), (63916,0.058079), (63917,0.060460), (63918,-0.134571), (63919,-0.204649), (63920,-0.336049), (63921,-0.048931), (63922,0.242364), (63923,0.179248), (63924,0.021844), (63925,0.167285), (63926,0.099986), (63927,0.065674), (63928,0.020210), (63929,-0.094465), (63930,0.213555), (63931,0.039889), (63932,0.061775), (63933,-0.042211), (63934,-0.182433), (63935,-0.360276), (63936,-0.074560), (63937,-0.217562), (63938,0.114608), (63939,-0.022364), (63940,0.124474), (63941,-0.043149), (63942,-0.008258), (63943,-0.167058), (63944,-0.282196), (63945,0.001202), (63946,0.281815), (63947,0.203370), (63948,0.049216), (63949,0.067389), (63950,-0.126252), (63951,-0.177289), (63952,-0.292891), (63953,-0.019248), (63954,0.217239), (63955,0.154123), (63956,-0.004215), (63957,0.124508), (63958,0.076258), (63959,0.008965), (63960,0.206898), (63961,0.012331), (63962,-0.011305), (63963,0.207066), (63964,0.244744), (63965,0.108705), (63966,0.089721), (63967,-0.155478), (63968,0.130707), (63969,0.006746), (63970,-0.073558), (63971,0.147136), (63972,0.317199), (63973,0.155612), (63974,0.109684), (63975,0.020094), (63976,-0.044882), (63977,0.220865), (63978,0.080649), (63979,0.442081), (63980,0.297682), (63981,0.274046), (63982,0.109209), (63983,0.080463), (63984,-0.054180), (63985,0.205531), (63986,0.039298), (63987,0.372859), (63988,0.215454), (63989,0.366469), (63990,0.238325), (63991,0.227701), (63992,0.383361), (63993,0.222707), (63994,0.240874), (63995,0.425338), (63996,0.438402), (63997,0.266132), (63998,0.216949), (63999,0.064191), (64000,0.365704), (64001,0.244993), (64002,0.203242), (64003,0.416504), (64004,0.579597), (64005,0.421723), (64006,0.323774), (64007,0.309430), (64008,0.090248), (64009,0.326734), (64010,0.154458), (64011,0.485239), (64012,0.364528), (64013,0.347861), (64014,0.198353), (64015,0.107830), (64016,-0.036106), (64017,0.292815), (64018,0.103358), (64019,0.489410), (64020,0.305525), (64021,0.462582), (64022,0.318177), (64023,0.361898), (64024,0.308074), (64025,0.183180), (64026,0.110315), (64027,0.296633), (64028,0.296691), (64029,0.147176), (64030,0.153277), (64031,-0.053833), (64032,0.202159), (64033,0.054973), (64034,0.055495), (64035,0.258068), (64036,0.403046), (64037,0.258647), (64038,0.187635), (64039,0.165395), (64040,0.394912), (64041,0.220783), (64042,0.180898), (64043,0.435030), (64044,0.453666), (64045,0.224729), (64046,0.167655), (64047,0.013031), (64048,0.312691), (64049,0.177579), (64050,0.114926), (64051,0.309609), (64052,0.447155), (64053,0.322724), (64054,0.282839), (64055,0.193249), (64056,0.350306), (64057,0.205437), (64058,0.191094), (64059,0.409928), (64060,0.398841), (64061,0.279520), (64062,0.225696), (64063,0.059463), (64064,0.316851), (64065,0.154800), (64066,0.129304), (64067,0.334207), (64068,0.511702), (64069,0.399813), (64070,0.344130), (64071,0.248040), (64072,0.469192), (64073,0.314574), (64074,0.255641), (64075,0.499553), (64076,0.497288), (64077,0.340347), (64078,0.229855), (64079,0.084987), (64080,0.384178), (64081,0.217018), (64082,0.196174), (64083,0.440093), (64084,0.581352), (64085,0.420698), (64086,0.345040), (64087,0.300972), (64088,0.399037), (64089,0.237914), (64090,0.189663), (64091,0.405705), (64092,0.439206), (64093,0.272973), (64094,0.266068), (64095,0.089616), (64096,0.383234), (64097,0.157546), (64098,0.131587), (64099,0.314654), (64100,0.461492), (64101,0.339855), (64102,0.285098), (64103,0.230348), (64104,0.359071), (64105,0.239286), (64106,0.586316), (64107,0.437271), (64108,0.433616), (64109,0.257627), (64110,0.174073), (64111,0.037107), (64112,0.350700), (64113,0.164955), (64114,0.467395), (64115,0.324856), (64116,0.477267), (64117,0.297102), (64118,0.360327), (64119,0.228934), (64120,0.251284), (64121,0.092483), (64122,0.472036), (64123,0.329954), (64124,0.286813), (64125,0.165639), (64126,0.072329), (64127,-0.048845), (64128,0.155124), (64129,0.000043), (64130,0.319202), (64131,0.179449), (64132,0.251967), (64133,0.153085), (64134,0.162898), (64135,0.033822), (64136,-0.120796), (64137,0.181181), (64138,0.419527), (64139,0.355948), (64140,0.204110), (64141,0.220893), (64142,0.052337), (64143,0.013842), (64144,-0.151465), (64145,0.123575), (64146,0.321508), (64147,0.282543), (64148,0.157656), (64149,0.326785), (64150,0.261352), (64151,0.233540), (64152,-0.143111), (64153,0.097552), (64154,0.303844), (64155,0.288110), (64156,0.139065), (64157,0.124722), (64158,-0.041512), (64159,-0.089762), (64160,-0.289903), (64161,-0.056203), (64162,0.210934), (64163,0.133886), (64164,0.045222), (64165,0.207389), (64166,0.147992), (64167,0.079767), (64168,-0.143135), (64169,0.125869), (64170,0.363282), (64171,0.296452), (64172,0.165986), (64173,0.167897), (64174,-0.027597), (64175,-0.073524), (64176,-0.224429), (64177,0.019020), (64178,0.280127), (64179,0.260674), (64180,0.062394), (64181,0.282618), (64182,0.135896), (64183,0.076030), (64184,-0.252312), (64185,-0.006533), (64186,0.272220), (64187,0.236048), (64188,0.042407), (64189,0.058720), (64190,-0.103793), (64191,-0.165513), (64192,-0.300162), (64193,-0.059963), (64194,0.184419), (64195,0.145461), (64196,-0.009627), (64197,0.187843), (64198,0.094997), (64199,0.023991), (64200,-0.157107), (64201,0.088665), (64202,0.318182), (64203,0.310807), (64204,0.182664), (64205,0.185045), (64206,0.051792), (64207,-0.017360), (64208,-0.195672), (64209,0.079830), (64210,0.340005), (64211,0.333557), (64212,0.159427), (64213,0.332276), (64214,0.246405), (64215,0.157742), (64216,-0.276504), (64217,-0.007037), (64218,0.277288), (64219,0.236934), (64220,0.099034), (64221,0.092587), (64222,-0.108480), (64223,-0.184139), (64224,-0.371267), (64225,-0.100880), (64226,0.215036), (64227,0.155176), (64228,-0.003625), (64229,0.145999), (64230,0.065232), (64231,0.014195), (64232,-0.154825), (64233,0.105812), (64234,0.403143), (64235,0.341424), (64236,0.162648), (64237,0.168279), (64238,-0.013746), (64239,-0.033193), (64240,-0.211968), (64241,0.095582), (64242,0.330671), (64243,0.251770), (64244,0.091573), (64245,0.273251), (64246,0.139065), (64247,0.117288), (64248,0.062074), (64249,0.330608), (64250,0.230799), (64251,0.530916), (64252,0.376298), (64253,0.389825), (64254,0.273760), (64255,0.219004), (64256,0.002145), (64257,0.307372), (64258,0.170869), (64259,0.515582), (64260,0.327984), (64261,0.474352), (64262,0.328557), (64263,0.405721), (64264,0.066234), (64265,0.364961), (64266,0.209874), (64267,0.560623), (64268,0.432016), (64269,0.440897), (64270,0.244013), (64271,0.130728), (64272,-0.010421), (64273,0.281807), (64274,0.108604), (64275,0.505803), (64276,0.319601), (64277,0.418593), (64278,0.296956), (64279,0.330451), (64280,0.425267), (64281,0.259497), (64282,0.168517), (64283,0.380845), (64284,0.428279), (64285,0.302922), (64286,0.259318), (64287,0.045245), (64288,0.334217), (64289,0.175416), (64290,0.145280), (64291,0.375261), (64292,0.526282), (64293,0.350756), (64294,0.296006), (64295,0.216634), (64296,0.193931), (64297,0.061605), (64298,0.390989), (64299,0.238688), (64300,0.276373), (64301,0.121749), (64302,0.003361), (64303,-0.090876), (64304,0.168372), (64305,0.027223), (64306,0.367753), (64307,0.218245), (64308,0.290763), (64309,0.163546), (64310,0.181256), (64311,0.042893), (64312,0.367162), (64313,0.206044), (64314,0.144318), (64315,0.409602), (64316,0.405947), (64317,0.230885), (64318,0.195176), (64319,0.031266), (64320,0.289117), (64321,0.155401), (64322,0.104827), (64323,0.335277), (64324,0.481182), (64325,0.343752), (64326,0.273667), (64327,0.216124), (64328,0.423813), (64329,0.236215), (64330,0.193537), (64331,0.450924), (64332,0.488603), (64333,0.318193), (64334,0.256937), (64335,0.081881), (64336,0.339262), (64337,0.208332), (64338,0.148009), (64339,0.354301), (64340,0.550838), (64341,0.363703), (64342,0.308483), (64343,0.236081), (64344,0.434478), (64345,0.257099), (64346,0.207915), (64347,0.456010), (64348,0.464428), (64349,0.329321), (64350,0.320087), (64351,0.091149), (64352,0.394986), (64353,0.218997), (64354,0.147985), (64355,0.375643), (64356,0.522017), (64357,0.327450), (64358,0.284772), (64359,0.225375), (64360,0.301613), (64361,0.184615), (64362,0.527932), (64363,0.381673), (64364,0.416565), (64365,0.245229), (64366,0.173753), (64367,-0.012918), (64368,0.247256), (64369,0.091705), (64370,0.466612), (64371,0.331499), (64372,0.464862), (64373,0.349724), (64374,0.329344), (64375,0.184945), (64376,0.202655), (64377,0.022483), (64378,0.408072), (64379,0.265064), (64380,0.292529), (64381,0.145801), (64382,0.005585), (64383,-0.130924), (64384,-0.319912), (64385,0.030374), (64386,-0.133073), (64387,0.208854), (64388,0.082100), (64389,0.256345), (64390,0.087326), (64391,0.120358), (64392,-0.141097), (64393,0.095389), (64394,-0.044833), (64395,0.290594), (64396,0.156872), (64397,0.126272), (64398,-0.023699), (64399,-0.099357), (64400,-0.246079), (64401,0.046142), (64402,-0.115445), (64403,0.228805), (64404,0.059322), (64405,0.192684), (64406,0.068260), (64407,0.075751), (64408,-0.036137), (64409,-0.221412), (64410,0.072206), (64411,0.310082), (64412,0.211663), (64413,0.113713), (64414,0.122130), (64415,-0.104021), (64416,-0.140662), (64417,-0.288311), (64418,-0.002589), (64419,0.216245), (64420,0.184250), (64421,0.039381), (64422,0.182043), (64423,0.070618), (64424,-0.254004), (64425,-0.423487), (64426,0.242187), (64427,0.090355), (64428,0.046287), (64429,-0.068387), (64430,-0.079018), (64431,-0.225740), (64432,-0.277241), (64433,-0.404921), (64434,0.264473), (64435,0.105672), (64436,0.062067), (64437,-0.116708), (64438,0.114669), (64439,-0.041809), (64440,-0.035715), (64441,-0.242361), (64442,0.019210), (64443,0.281244), (64444,0.204189), (64445,0.074656), (64446,0.089109), (64447,-0.093843), (64448,-0.156025), (64449,-0.310650), (64450,-0.020282), (64451,0.234320), (64452,0.178636), (64453,-0.033583), (64454,0.141589), (64455,0.078010), (64456,0.024186), (64457,-0.146230), (64458,0.121377), (64459,0.408495), (64460,0.344446), (64461,0.154525), (64462,0.168521), (64463,0.014830), (64464,-0.073370), (64465,-0.182465), (64466,0.085135), (64467,0.348565), (64468,0.294735), (64469,0.107601), (64470,0.263268), (64471,0.189469), (64472,-0.019963), (64473,-0.173191), (64474,0.126933), (64475,0.374565), (64476,0.271036), (64477,0.171226), (64478,0.143883), (64479,-0.033032), (64480,-0.091972), (64481,-0.235907), (64482,0.061893), (64483,0.321604), (64484,0.238513), (64485,0.080639), (64486,0.254885), (64487,0.170404), (64488,0.111934), (64489,-0.072414), (64490,0.182187), (64491,0.446538), (64492,0.382495), (64493,0.182355), (64494,0.232112), (64495,0.085390), (64496,0.058041), (64497,-0.129094), (64498,0.171956), (64499,0.403333), (64500,0.313279), (64501,0.166551), (64502,0.306889), (64503,0.236341), (64504,0.092869), (64505,-0.064999), (64506,0.180774), (64507,0.487397), (64508,0.421494), (64509,0.249688), (64510,0.285050), (64511,0.112310), (64512,-0.023729), (64513,-0.189029), (64514,0.069749), (64515,0.346641), (64516,0.303500), (64517,0.143309), (64518,0.325914), (64519,0.213562), (64520,-0.008412), (64521,-0.194151), (64522,0.128265), (64523,0.304363), (64524,0.294666), (64525,0.113574), (64526,0.146142), (64527,-0.019628), (64528,-0.064159), (64529,-0.232252), (64530,0.078091), (64531,0.340588), (64532,0.222657), (64533,0.072686), (64534,0.208378), (64535,0.161054), (64536,-0.112010), (64537,0.154664), (64538,0.040452), (64539,0.358228), (64540,0.226365), (64541,0.248721), (64542,0.053220), (64543,-0.025681), (64544,-0.127814), (64545,0.113776), (64546,-0.049201), (64547,0.269494), (64548,0.151570), (64549,0.302591), (64550,0.154472), (64551,0.172182), (64552,-0.033068), (64553,0.307463), (64554,0.109182), (64555,0.482693), (64556,0.331325), (64557,0.344382), (64558,0.223208), (64559,0.115966), (64560,-0.021470), (64561,0.205730), (64562,0.065044), (64563,0.400928), (64564,0.249560), (64565,0.461426), (64566,0.239921), (64567,0.219071), (64568,-0.150604), (64569,0.197822), (64570,0.047381), (64571,0.335426), (64572,0.226324), (64573,0.286770), (64574,0.130286), (64575,0.017008), (64576,-0.127854), (64577,0.151361), (64578,-0.032060), (64579,0.287575), (64580,0.174754), (64581,0.333207), (64582,0.230611), (64583,0.208835), (64584,-0.081881), (64585,0.193159), (64586,0.032035), (64587,0.372102), (64588,0.191004), (64589,0.234724), (64590,0.069418), (64591,0.025813), (64592,-0.113940), (64593,0.116968), (64594,-0.019535), (64595,0.301484), (64596,0.206320), (64597,0.356878), (64598,0.207826), (64599,0.213457), (64600,-0.018267), (64601,0.234475), (64602,0.085430), (64603,0.411565), (64604,0.246721), (64605,0.252816), (64606,0.088906), (64607,0.063879), (64608,-0.103744), (64609,0.140638), (64610,0.000416), (64611,0.344202), (64612,0.201657), (64613,0.349422), (64614,0.246826), (64615,0.230159), (64616,-0.127907), (64617,0.119725), (64618,0.411483), (64619,0.363232), (64620,0.207218), (64621,0.206349), (64622,0.024324), (64623,-0.013708), (64624,-0.159503), (64625,0.120646), (64626,0.360382), (64627,0.306089), (64628,0.162154), (64629,0.271835), (64630,0.214292), (64631,0.148852), (64632,-0.042922), (64633,0.226538), (64634,0.122546), (64635,0.401768), (64636,0.267119), (64637,0.289938), (64638,0.095834), (64639,0.034578), (64640,-0.304910), (64641,-0.061924), (64642,-0.207256), (64643,0.143030), (64644,-0.010191), (64645,0.111099), (64646,-0.034233), (64647,-0.007237), (64648,-0.252430), (64649,0.033286), (64650,-0.150130), (64651,0.202479), (64652,0.065977), (64653,0.092509), (64654,-0.039817), (64655,-0.155882), (64656,-0.305860), (64657,-0.016888), (64658,-0.178475), (64659,0.175060), (64660,0.024625), (64661,0.195151), (64662,0.016839), (64663,0.041518), (64664,-0.097314), (64665,-0.270047), (64666,0.006382), (64667,0.287928), (64668,0.244317), (64669,0.067871), (64670,0.094403), (64671,-0.125712), (64672,-0.181395), (64673,-0.315575), (64674,-0.042865), (64675,0.208950), (64676,0.135152), (64677,-0.027826), (64678,0.138517), (64679,0.073548), (64680,-0.265946), (64681,-0.434496), (64682,0.305961), (64683,0.123009), (64684,0.106806), (64685,-0.050135), (64686,-0.099776), (64687,-0.246968), (64688,-0.316583), (64689,-0.446123), (64690,0.257184), (64691,0.092340), (64692,0.051986), (64693,-0.078944), (64694,0.151036), (64695,-0.030056), (64696,-0.127079), (64697,-0.286806), (64698,0.008665), (64699,0.267912), (64700,0.225234), (64701,0.073403), (64702,0.087856), (64703,-0.123429), (64704,-0.175863), (64705,-0.353705), (64706,-0.024791), (64707,0.199623), (64708,0.134184), (64709,-0.004642), (64710,0.126398), (64711,0.092549), (64712,0.001562), (64713,-0.199968), (64714,0.048591), (64715,0.320380), (64716,0.286525), (64717,0.123548), (64718,0.105021), (64719,-0.067248), (64720,-0.095988), (64721,-0.274763), (64722,0.026287), (64723,0.260914), (64724,0.219163), (64725,0.110067), (64726,0.223925), (64727,0.173351), (64728,-0.060696), (64729,-0.215784), (64730,0.089450), (64731,0.303638), (64732,0.243772), (64733,0.106806), (64734,0.154240), (64735,-0.007811), (64736,-0.055598), (64737,-0.252952), (64738,0.028587), (64739,0.246958), (64740,0.182915), (64741,0.002750), (64742,0.161660), (64743,0.116659), (64744,0.047507), (64745,-0.132658), (64746,0.180934), (64747,0.370502), (64748,0.319001), (64749,0.187145), (64750,0.189056), (64751,0.000995), (64752,-0.040757), (64753,-0.181906), (64754,0.114499), (64755,0.333797), (64756,0.282759), (64757,0.102131), (64758,0.257328), (64759,0.201644), (64760,0.009864), (64761,-0.144291), (64762,0.142821), (64763,0.340291), (64764,0.325947), (64765,0.193157), (64766,0.237341), (64767,0.008404), (64768,-0.059822), (64769,-0.198648), (64770,0.098689), (64771,0.324024), (64772,0.272523), (64773,0.128118), (64774,0.254054), (64775,0.170500), (64776,-0.037536), (64777,-0.191227), (64778,0.070344), (64779,0.322622), (64780,0.280407), (64781,0.114637), (64782,0.156035), (64783,-0.063147), (64784,-0.086783), (64785,-0.233505), (64786,0.022956), (64787,0.293813), (64788,0.207472), (64789,0.064000), (64790,0.185290), (64791,0.150508), (64792,-0.000860), (64793,0.291831), (64794,0.149749), (64795,0.110328), (64796,0.317083), (64797,0.377059), (64798,0.205717), (64799,0.116126), (64800,-0.064972), (64801,0.209604), (64802,0.071241), (64803,0.033210), (64804,0.249258), (64805,0.401669), (64806,0.217784), (64807,0.189971), (64808,-0.083562), (64809,0.186368), (64810,0.070766), (64811,0.427088), (64812,0.294768), (64813,0.240012), (64814,0.077961), (64815,0.065477), (64816,-0.074282), (64817,0.199831), (64818,0.014086), (64819,0.346257), (64820,0.173988), (64821,0.331508), (64822,0.179213), (64823,0.178802), (64824,-0.116560), (64825,0.162662), (64826,-0.007290), (64827,0.303516), (64828,0.164220), (64829,0.207941), (64830,-0.003345), (64831,-0.072034), (64832,-0.203427), (64833,0.061387), (64834,-0.076976), (64835,0.283066), (64836,0.036013), (64837,0.204679), (64838,0.033806), (64839,0.120720), (64840,-0.153740), (64841,0.134768), (64842,0.005698), (64843,0.370849), (64844,0.217621), (64845,0.195382), (64846,0.028222), (64847,-0.053009), (64848,-0.167221), (64849,0.114788), (64850,-0.055628), (64851,0.263537), (64852,0.093591), (64853,0.233460), (64854,0.162911), (64855,0.143464), (64856,0.049691), (64857,0.323334), (64858,0.165460), (64859,0.119069), (64860,0.297960), (64861,0.376051), (64862,0.231183), (64863,0.157384), (64864,-0.007453), (64865,0.269910), (64866,0.150126), (64867,0.076327), (64868,0.292376), (64869,0.458718), (64870,0.317570), (64871,0.270245), (64872,-0.154244), (64873,0.121259), (64874,0.369817), (64875,0.326213), (64876,0.173918), (64877,0.160971), (64878,0.019352), (64879,-0.040045), (64880,-0.185376), (64881,0.064115), (64882,0.308961), (64883,0.250028), (64884,0.090764), (64885,0.221803), (64886,0.185168), (64887,0.111370), (64888,-0.046968), (64889,0.209493), (64890,0.062771), (64891,0.410265), (64892,0.260756), (64893,0.273357), (64894,0.105264), (64895,0.081170), (64896,-0.288511), (64897,0.007893), (64898,-0.193180), (64899,0.167325), (64900,-0.017950), (64901,0.114023), (64902,-0.036419), (64903,0.007302), (64904,-0.240214), (64905,0.034819), (64906,-0.102610), (64907,0.242103), (64908,0.064254), (64909,0.104262), (64910,-0.089379), (64911,-0.159928), (64912,-0.327551), (64913,-0.028824), (64914,-0.195520), (64915,0.197965), (64916,0.012684), (64917,0.101000), (64918,-0.027613), (64919,0.026790), (64920,0.027311), (64921,-0.188157), (64922,0.118466), (64923,0.014480), (64924,0.337822), (64925,0.191563), (64926,0.214846), (64927,0.060228), (64928,-0.032155), (64929,-0.176554), (64930,0.098486), (64931,-0.011079), (64932,0.313195), (64933,0.192015), (64934,0.244095), (64935,0.124317), (64936,-0.075823), (64937,-0.229051), (64938,0.084072), (64939,0.298260), (64940,0.238864), (64941,0.065198), (64942,0.094523), (64943,-0.087502), (64944,-0.112528), (64945,-0.257397), (64946,-0.034379), (64947,0.183522), (64948,0.165929), (64949,-0.021669), (64950,0.142351), (64951,0.071345), (64952,-0.199865), (64953,-0.363312), (64954,-0.044610), (64955,0.211381), (64956,0.116681), (64957,-0.083922), (64958,-0.057853), (64959,-0.262640), (64960,-0.299745), (64961,-0.419992), (64962,-0.141233), (64963,0.105466), (64964,0.043283), (64965,-0.121091), (64966,0.003449), (64967,-0.049448), (64968,-0.113490), (64969,-0.278790), (64970,0.052447), (64971,0.277318), (64972,0.233714), (64973,0.108820), (64974,0.093549), (64975,-0.080110), (64976,-0.146013), (64977,-0.324788), (64978,-0.032097), (64979,0.198810), (64980,0.146376), (64981,-0.054227), (64982,0.118158), (64983,0.034604), (64984,-0.045230), (64985,-0.183593), (64986,0.086337), (64987,-0.027874), (64988,0.327058), (64989,0.169184), (64990,0.164132), (64991,0.035062), (64992,-0.092618), (64993,-0.241663), (64994,0.056131), (64995,-0.106846), (64996,0.239257), (64997,0.158959), (64998,0.282573), (64999,0.091255), (65000,0.142409), (65001,0.015192), (65002,0.269330), (65003,0.140253), (65004,0.422725), (65005,0.234658), (65006,0.307176), (65007,0.140016), (65008,0.025811), (65009,-0.139959), (65010,0.202894), (65011,0.008790), (65012,0.405989), (65013,0.198422), (65014,0.388453), (65015,0.251487), (65016,0.198590), (65017,0.001236), (65018,0.289281), (65019,0.177856), (65020,0.503991), (65021,0.321966), (65022,0.359644), (65023,0.203630), (65024,0.143306), (65025,0.022595), (65026,0.299025), (65027,0.128609), (65028,0.438952), (65029,0.255993), (65030,0.457176), (65031,0.286303), (65032,0.155373), (65033,0.023047), (65034,0.272539), (65035,0.110019), (65036,0.465884), (65037,0.321479), (65038,0.274624), (65039,0.138585), (65040,0.071286), (65041,-0.046638), (65042,0.231187), (65043,0.023151), (65044,0.399912), (65045,0.226715), (65046,0.369370), (65047,0.241227), (65048,0.036441), (65049,0.340277), (65050,0.200519), (65051,0.140659), (65052,0.374352), (65053,0.381379), (65054,0.245340), (65055,0.139025), (65056,-0.025812), (65057,0.263623), (65058,0.092750), (65059,0.009659), (65060,0.236389), (65061,0.393910), (65062,0.247651), (65063,0.219839), (65064,-0.036043), (65065,0.260831), (65066,0.082055), (65067,0.069571), (65068,0.335318), (65069,0.326547), (65070,0.181685), (65071,0.133435), (65072,-0.075998), (65073,0.248740), (65074,0.098299), (65075,0.039366), (65076,0.283748), (65077,0.398069), (65078,0.237415), (65079,0.207743), (65080,0.014102), (65081,0.268240), (65082,0.139633), (65083,0.102528), (65084,0.348300), (65085,0.322811), (65086,0.182595), (65087,0.139454), (65088,-0.047681), (65089,0.269161), (65090,0.100142), (65091,0.054677), (65092,0.260037), (65093,0.450074), (65094,0.282451), (65095,0.184495), (65096,0.033590), (65097,0.305379), (65098,0.158658), (65099,0.141527), (65100,0.378477), (65101,0.411972), (65102,0.202083), (65103,0.138967), (65104,0.008037), (65105,0.245450), (65106,0.085722), (65107,0.066269), (65108,0.282781), (65109,0.400815), (65110,0.247593), (65111,0.228603), (65112,0.093027), (65113,0.354128), (65114,0.225058), (65115,0.175880), (65116,0.410507), (65117,0.437039), (65118,0.266623), (65119,0.236957), (65120,0.001050), (65121,0.265401), (65122,0.128898), (65123,0.069032), (65124,0.311091), (65125,0.440741), (65126,0.293092), (65127,0.236482), (65128,-0.024972), (65129,0.262139), (65130,0.116344), (65131,0.496361), (65132,0.326878), (65133,0.342728), (65134,0.204365), (65135,0.093867), (65136,-0.110450), (65137,0.140895), (65138,0.027154), (65139,0.335637), (65140,0.196341), (65141,0.374300), (65142,0.284709), (65143,0.305669), (65144,-0.161093), (65145,0.107910), (65146,-0.049964), (65147,0.315650), (65148,0.223273), (65149,0.202430), (65150,0.068244), (65151,-0.064546), (65152,-0.091895), (65153,-0.227001), (65154,0.027600), (65155,0.207875), (65156,0.197251), (65157,0.056102), (65158,0.206189), (65159,0.101734), (65160,-0.051024), (65161,-0.217721), (65162,0.074501), (65163,0.327242), (65164,0.235792), (65165,0.093253), (65166,0.069153), (65167,-0.081751), (65168,-0.110954), (65169,-0.263718), (65170,0.002955), (65171,0.239442), (65172,0.166107), (65173,0.017062), (65174,0.148571), (65175,0.121222), (65176,-0.050115), (65177,-0.195910), (65178,0.107457), (65179,0.366241), (65180,0.294303), (65181,0.151294), (65182,0.163888), (65183,-0.050185), (65184,-0.093789), (65185,-0.249803), (65186,0.018730), (65187,0.255216), (65188,0.237623), (65189,0.068603), (65190,0.231696), (65191,0.164404), (65192,-0.151865), (65193,-0.227981), (65194,0.021041), (65195,0.288648), (65196,0.114056), (65197,0.043507), (65198,-0.051193), (65199,-0.109193), (65200,-0.235946), (65201,-0.295806), (65202,-0.064899), (65203,0.212000), (65204,0.062022), (65205,0.020277), (65206,-0.080002), (65207,0.128614), (65208,-0.085922), (65209,-0.134643), (65210,-0.274859), (65211,0.389425), (65212,0.231088), (65213,0.165649), (65214,-0.008480), (65215,0.002260), (65216,-0.173723), (65217,-0.228479), (65218,-0.346867), (65219,0.305808), (65220,0.153043), (65221,0.107579), (65222,-0.071660), (65223,0.166216), (65224,-0.010699), (65225,-0.034329), (65226,-0.230286), (65227,0.499488), (65228,0.316536), (65229,0.263176), (65230,0.090906), (65231,0.091891), (65232,-0.106859), (65233,-0.133275), (65234,-0.229835), (65235,0.420047), (65236,0.251960), (65237,0.135426), (65238,-0.021052), (65239,0.222404), (65240,-0.089682), (65241,-0.145829), (65242,-0.308343), (65243,0.374056), (65244,0.217115), (65245,0.160968), (65246,0.019813), (65247,0.031023), (65248,-0.170050), (65249,-0.170456), (65250,-0.358054), (65251,0.250025), (65252,0.105157), (65253,0.105215), (65254,-0.047080), (65255,0.166645), (65256,0.020387), (65257,-0.029260), (65258,-0.178305), (65259,0.482729), (65260,0.322532), (65261,0.263135), (65262,0.143814), (65263,0.109502), (65264,-0.069273), (65265,-0.073861), (65266,-0.217334), (65267,0.449273), (65268,0.296972), (65269,0.273342), (65270,0.103859), (65271,0.346382), (65272,0.041728), (65273,-0.010699), (65274,-0.189938), (65275,0.473419), (65276,0.351312), (65277,0.265898), (65278,0.122426), (65279,0.122947), (65280,-0.019592), (65281,-0.074812), (65282,-0.217357), (65283,0.435781), (65284,0.272334), (65285,0.229193), (65286,0.096410), (65287,0.274831), (65288,-0.052584), (65289,-0.097578), (65290,-0.249416), (65291,0.458994), (65292,0.314595), (65293,0.277490), (65294,0.087105), (65295,0.047684), (65296,-0.097185), (65297,-0.166337), (65298,-0.307486), (65299,0.398137), (65300,0.225868), (65301,0.156252), (65302,0.022999), (65303,0.231608), (65304,0.095569), (65305,-0.067408), (65306,0.198339), (65307,0.072519), (65308,0.436737), (65309,0.333677), (65310,0.307725), (65311,0.136845), (65312,0.089058), (65313,-0.065560), (65314,0.183932), (65315,0.012126), (65316,0.404214), (65317,0.257956), (65318,0.343016), (65319,0.206044), (65320,0.049103), (65321,-0.105985), (65322,0.175561), (65323,0.441308), (65324,0.387014), (65325,0.153430), (65326,0.179499), (65327,0.017449), (65328,0.005892), (65329,-0.165914), (65330,0.136996), (65331,0.373482), (65332,0.326158), (65333,0.158065), (65334,0.330450), (65335,0.252006), (65336,0.022605), (65337,-0.165457), (65338,0.108650), (65339,0.322838), (65340,0.303385), (65341,0.152480), (65342,0.188305), (65343,-0.031810), (65344,-0.082847), (65345,-0.236538), (65346,-0.002839), (65347,0.251763), (65348,0.222090), (65349,0.043315), (65350,0.190153), (65351,0.094526), (65352,-0.052665), (65353,-0.181272), (65354,0.140216), (65355,0.303310), (65356,0.311727), (65357,0.120409), (65358,0.172959), (65359,-0.039260), (65360,-0.033629), (65361,-0.198002), (65362,0.064495), (65363,0.274500), (65364,0.278272), (65365,0.125050), (65366,0.250980), (65367,0.132593), (65368,0.160058), (65369,0.009153), (65370,0.282796), (65371,0.129105), (65372,0.474745), (65373,0.342888), (65374,0.366165), (65375,0.188786), (65376,0.156327), (65377,-0.014083), (65378,0.255377), (65379,0.086827), (65380,0.474733), (65381,0.267630), (65382,0.464630), (65383,0.238942), (65384,-0.061992), (65385,-0.223579), (65386,0.475075), (65387,0.362723), (65388,0.238763), (65389,0.125015), (65390,0.063295), (65391,-0.063922), (65392,-0.169767), (65393,-0.297911), (65394,0.409572), (65395,0.194104), (65396,0.163968), (65397,0.032105), (65398,0.295066), (65399,0.129302), (65400,0.026243), (65401,-0.098188), (65402,0.163377), (65403,0.408692), (65404,0.334424), (65405,0.191421), (65406,0.173828), (65407,0.015954), (65408,-0.153529), (65409,-0.303970), (65410,0.002653), (65411,0.264223), (65412,0.200181), (65413,0.031624), (65414,0.208186), (65415,0.139497), (65416,-0.003511), (65417,-0.176244), (65418,0.102045), (65419,0.292082), (65420,0.247545), (65421,0.068776), (65422,0.079510), (65423,-0.113198), (65424,-0.119176), (65425,-0.269154), (65426,-0.008047), (65427,0.209391), (65428,0.167640), (65429,0.031601), (65430,0.184012), (65431,0.100464), (65432,-0.070416), (65433,-0.111697), (65434,-0.299295), (65435,0.383567), (65436,0.265642), (65437,0.240616), (65438,0.040939), (65439,0.036351), (65440,-0.071817), (65441,-0.111246), (65442,-0.277479), (65443,0.370550), (65444,0.223364), (65445,0.159785), (65446,0.025136), (65447,0.237001), (65448,-0.176806), (65449,-0.229703), (65450,-0.012259), (65451,0.293432), (65452,0.115126), (65453,0.062229), (65454,-0.125832), (65455,-0.135530), (65456,-0.285971), (65457,-0.291486), (65458,-0.044787), (65459,0.251617), (65460,0.100249), (65461,0.034346), (65462,-0.058030), (65463,0.132470), (65464,-0.063950), (65465,-0.134962), (65466,-0.284477), (65467,0.404428), (65468,0.256773), (65469,0.183444), (65470,0.012101), (65471,-0.011535), (65472,-0.118771), (65473,-0.153553), (65474,-0.280769), (65475,0.349144), (65476,0.184301), (65477,0.106326), (65478,-0.030647), (65479,0.192834), (65480,-0.075120), (65481,-0.112688), (65482,-0.221327), (65483,0.436458), (65484,0.292059), (65485,0.260527), (65486,0.106372), (65487,0.072987), (65488,-0.097893), (65489,-0.171228), (65490,-0.295188), (65491,0.374668), (65492,0.171278), (65493,0.161117), (65494,0.039010), (65495,0.281996), (65496,0.048875), (65497,-0.039319), (65498,-0.213448), (65499,0.446653), (65500,0.270207), (65501,0.188043), (65502,0.053400), (65503,0.049739), (65504,-0.085838), (65505,-0.102498), (65506,-0.258976), (65507,0.448038), (65508,0.250684), (65509,0.181995), (65510,0.033883), (65511,0.282442), (65512,-0.120220), (65513,-0.175903), (65514,-0.283145), (65515,0.389041), (65516,0.197260), (65517,0.186629), (65518,0.034798), (65519,-0.044110), (65520,-0.217769), (65521,-0.288318), (65522,-0.404852), (65523,0.331428), (65524,0.185639), (65525,0.099762), (65526,-0.031631), (65527,0.199276), (65528,-0.075647), (65529,-0.089058), (65530,-0.252968), (65531,0.411779), (65532,0.219998), (65533,0.172680), (65534,-0.020034), (65535,-0.000001), 
.ends AD3552R_INL